-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 13 2021 17:23:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zim" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zim
entity zim is
port (
    VAC_DRDY : in std_logic;
    IAC_FLT1 : out std_logic;
    DDS_SCK : out std_logic;
    ICE_IOR_166 : in std_logic;
    ICE_IOR_119 : in std_logic;
    DDS_MOSI : out std_logic;
    VAC_MISO : in std_logic;
    DDS_MOSI1 : out std_logic;
    ICE_IOR_146 : in std_logic;
    VDC_CLK : out std_logic;
    ICE_IOT_222 : in std_logic;
    IAC_CS : out std_logic;
    ICE_IOL_18B : in std_logic;
    ICE_IOL_13A : in std_logic;
    ICE_IOB_81 : in std_logic;
    VAC_OSR1 : out std_logic;
    IAC_MOSI : out std_logic;
    DDS_CS1 : out std_logic;
    ICE_IOL_4B : in std_logic;
    ICE_IOB_94 : in std_logic;
    VAC_CS : out std_logic;
    VAC_CLK : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    ICE_IOR_167 : in std_logic;
    ICE_IOR_118 : in std_logic;
    RTD_SDO : in std_logic;
    IAC_OSR0 : out std_logic;
    VDC_SCLK : out std_logic;
    VAC_FLT1 : out std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_IOR_165 : in std_logic;
    ICE_IOR_147 : in std_logic;
    ICE_IOL_14A : in std_logic;
    ICE_IOL_13B : in std_logic;
    ICE_IOB_91 : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_RNG_0 : out std_logic;
    VDC_RNG0 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    ICE_IOR_152 : in std_logic;
    ICE_IOL_12A : in std_logic;
    RTD_DRDY : in std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_IOT_177 : in std_logic;
    ICE_IOR_141 : in std_logic;
    ICE_IOB_80 : in std_logic;
    ICE_IOB_102 : in std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    IAC_MISO : in std_logic;
    VAC_OSR0 : out std_logic;
    VAC_MOSI : out std_logic;
    TEST_LED : out std_logic;
    ICE_IOR_148 : in std_logic;
    STAT_COMM : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_IOR_161 : in std_logic;
    ICE_IOB_95 : in std_logic;
    ICE_IOB_82 : in std_logic;
    ICE_IOB_104 : in std_logic;
    IAC_CLK : out std_logic;
    DDS_CS : out std_logic;
    SELIRNG0 : out std_logic;
    RTD_SDI : out std_logic;
    ICE_IOT_221 : in std_logic;
    ICE_IOT_197 : in std_logic;
    DDS_MCLK : out std_logic;
    RTD_SCLK : out std_logic;
    RTD_CS : out std_logic;
    ICE_IOR_137 : in std_logic;
    IAC_OSR1 : out std_logic;
    VAC_FLT0 : out std_logic;
    ICE_IOR_144 : in std_logic;
    ICE_IOR_128 : in std_logic;
    ICE_GPMO_1 : in std_logic;
    IAC_SCLK : out std_logic;
    EIS_SYNCCLK : in std_logic;
    ICE_IOR_139 : in std_logic;
    ICE_IOL_4A : in std_logic;
    VAC_SCLK : out std_logic;
    THERMOSTAT : in std_logic;
    ICE_IOR_164 : in std_logic;
    ICE_IOB_103 : in std_logic;
    AMPV_POW : out std_logic;
    VDC_SDO : in std_logic;
    ICE_IOT_174 : in std_logic;
    ICE_IOR_140 : in std_logic;
    ICE_IOB_96 : in std_logic;
    CONT_SD : out std_logic;
    AC_ADC_SYNC : out std_logic;
    SELIRNG1 : out std_logic;
    ICE_IOL_12B : in std_logic;
    ICE_IOR_160 : in std_logic;
    ICE_IOR_136 : in std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_IOT_198 : in std_logic;
    ICE_IOT_173 : in std_logic;
    IAC_DRDY : in std_logic;
    ICE_IOT_178 : in std_logic;
    ICE_IOR_138 : in std_logic;
    ICE_IOR_120 : in std_logic;
    IAC_FLT0 : out std_logic;
    DDS_SCK1 : out std_logic);
end zim;

-- Architecture of zim
-- View name is \INTERFACE\
architecture \INTERFACE\ of zim is

signal \N__65921\ : std_logic;
signal \N__65920\ : std_logic;
signal \N__65919\ : std_logic;
signal \N__65912\ : std_logic;
signal \N__65911\ : std_logic;
signal \N__65910\ : std_logic;
signal \N__65903\ : std_logic;
signal \N__65902\ : std_logic;
signal \N__65901\ : std_logic;
signal \N__65894\ : std_logic;
signal \N__65893\ : std_logic;
signal \N__65892\ : std_logic;
signal \N__65885\ : std_logic;
signal \N__65884\ : std_logic;
signal \N__65883\ : std_logic;
signal \N__65876\ : std_logic;
signal \N__65875\ : std_logic;
signal \N__65874\ : std_logic;
signal \N__65867\ : std_logic;
signal \N__65866\ : std_logic;
signal \N__65865\ : std_logic;
signal \N__65858\ : std_logic;
signal \N__65857\ : std_logic;
signal \N__65856\ : std_logic;
signal \N__65849\ : std_logic;
signal \N__65848\ : std_logic;
signal \N__65847\ : std_logic;
signal \N__65840\ : std_logic;
signal \N__65839\ : std_logic;
signal \N__65838\ : std_logic;
signal \N__65831\ : std_logic;
signal \N__65830\ : std_logic;
signal \N__65829\ : std_logic;
signal \N__65822\ : std_logic;
signal \N__65821\ : std_logic;
signal \N__65820\ : std_logic;
signal \N__65813\ : std_logic;
signal \N__65812\ : std_logic;
signal \N__65811\ : std_logic;
signal \N__65804\ : std_logic;
signal \N__65803\ : std_logic;
signal \N__65802\ : std_logic;
signal \N__65795\ : std_logic;
signal \N__65794\ : std_logic;
signal \N__65793\ : std_logic;
signal \N__65786\ : std_logic;
signal \N__65785\ : std_logic;
signal \N__65784\ : std_logic;
signal \N__65777\ : std_logic;
signal \N__65776\ : std_logic;
signal \N__65775\ : std_logic;
signal \N__65768\ : std_logic;
signal \N__65767\ : std_logic;
signal \N__65766\ : std_logic;
signal \N__65759\ : std_logic;
signal \N__65758\ : std_logic;
signal \N__65757\ : std_logic;
signal \N__65750\ : std_logic;
signal \N__65749\ : std_logic;
signal \N__65748\ : std_logic;
signal \N__65741\ : std_logic;
signal \N__65740\ : std_logic;
signal \N__65739\ : std_logic;
signal \N__65732\ : std_logic;
signal \N__65731\ : std_logic;
signal \N__65730\ : std_logic;
signal \N__65723\ : std_logic;
signal \N__65722\ : std_logic;
signal \N__65721\ : std_logic;
signal \N__65714\ : std_logic;
signal \N__65713\ : std_logic;
signal \N__65712\ : std_logic;
signal \N__65705\ : std_logic;
signal \N__65704\ : std_logic;
signal \N__65703\ : std_logic;
signal \N__65696\ : std_logic;
signal \N__65695\ : std_logic;
signal \N__65694\ : std_logic;
signal \N__65687\ : std_logic;
signal \N__65686\ : std_logic;
signal \N__65685\ : std_logic;
signal \N__65678\ : std_logic;
signal \N__65677\ : std_logic;
signal \N__65676\ : std_logic;
signal \N__65669\ : std_logic;
signal \N__65668\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65660\ : std_logic;
signal \N__65659\ : std_logic;
signal \N__65658\ : std_logic;
signal \N__65651\ : std_logic;
signal \N__65650\ : std_logic;
signal \N__65649\ : std_logic;
signal \N__65642\ : std_logic;
signal \N__65641\ : std_logic;
signal \N__65640\ : std_logic;
signal \N__65633\ : std_logic;
signal \N__65632\ : std_logic;
signal \N__65631\ : std_logic;
signal \N__65624\ : std_logic;
signal \N__65623\ : std_logic;
signal \N__65622\ : std_logic;
signal \N__65615\ : std_logic;
signal \N__65614\ : std_logic;
signal \N__65613\ : std_logic;
signal \N__65606\ : std_logic;
signal \N__65605\ : std_logic;
signal \N__65604\ : std_logic;
signal \N__65597\ : std_logic;
signal \N__65596\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65588\ : std_logic;
signal \N__65587\ : std_logic;
signal \N__65586\ : std_logic;
signal \N__65579\ : std_logic;
signal \N__65578\ : std_logic;
signal \N__65577\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65569\ : std_logic;
signal \N__65568\ : std_logic;
signal \N__65561\ : std_logic;
signal \N__65560\ : std_logic;
signal \N__65559\ : std_logic;
signal \N__65552\ : std_logic;
signal \N__65551\ : std_logic;
signal \N__65550\ : std_logic;
signal \N__65543\ : std_logic;
signal \N__65542\ : std_logic;
signal \N__65541\ : std_logic;
signal \N__65534\ : std_logic;
signal \N__65533\ : std_logic;
signal \N__65532\ : std_logic;
signal \N__65525\ : std_logic;
signal \N__65524\ : std_logic;
signal \N__65523\ : std_logic;
signal \N__65516\ : std_logic;
signal \N__65515\ : std_logic;
signal \N__65514\ : std_logic;
signal \N__65507\ : std_logic;
signal \N__65506\ : std_logic;
signal \N__65505\ : std_logic;
signal \N__65498\ : std_logic;
signal \N__65497\ : std_logic;
signal \N__65496\ : std_logic;
signal \N__65489\ : std_logic;
signal \N__65488\ : std_logic;
signal \N__65487\ : std_logic;
signal \N__65480\ : std_logic;
signal \N__65479\ : std_logic;
signal \N__65478\ : std_logic;
signal \N__65471\ : std_logic;
signal \N__65470\ : std_logic;
signal \N__65469\ : std_logic;
signal \N__65462\ : std_logic;
signal \N__65461\ : std_logic;
signal \N__65460\ : std_logic;
signal \N__65453\ : std_logic;
signal \N__65452\ : std_logic;
signal \N__65451\ : std_logic;
signal \N__65444\ : std_logic;
signal \N__65443\ : std_logic;
signal \N__65442\ : std_logic;
signal \N__65435\ : std_logic;
signal \N__65434\ : std_logic;
signal \N__65433\ : std_logic;
signal \N__65426\ : std_logic;
signal \N__65425\ : std_logic;
signal \N__65424\ : std_logic;
signal \N__65417\ : std_logic;
signal \N__65416\ : std_logic;
signal \N__65415\ : std_logic;
signal \N__65408\ : std_logic;
signal \N__65407\ : std_logic;
signal \N__65406\ : std_logic;
signal \N__65399\ : std_logic;
signal \N__65398\ : std_logic;
signal \N__65397\ : std_logic;
signal \N__65390\ : std_logic;
signal \N__65389\ : std_logic;
signal \N__65388\ : std_logic;
signal \N__65381\ : std_logic;
signal \N__65380\ : std_logic;
signal \N__65379\ : std_logic;
signal \N__65372\ : std_logic;
signal \N__65371\ : std_logic;
signal \N__65370\ : std_logic;
signal \N__65363\ : std_logic;
signal \N__65362\ : std_logic;
signal \N__65361\ : std_logic;
signal \N__65354\ : std_logic;
signal \N__65353\ : std_logic;
signal \N__65352\ : std_logic;
signal \N__65345\ : std_logic;
signal \N__65344\ : std_logic;
signal \N__65343\ : std_logic;
signal \N__65336\ : std_logic;
signal \N__65335\ : std_logic;
signal \N__65334\ : std_logic;
signal \N__65327\ : std_logic;
signal \N__65326\ : std_logic;
signal \N__65325\ : std_logic;
signal \N__65318\ : std_logic;
signal \N__65317\ : std_logic;
signal \N__65316\ : std_logic;
signal \N__65309\ : std_logic;
signal \N__65308\ : std_logic;
signal \N__65307\ : std_logic;
signal \N__65300\ : std_logic;
signal \N__65299\ : std_logic;
signal \N__65298\ : std_logic;
signal \N__65291\ : std_logic;
signal \N__65290\ : std_logic;
signal \N__65289\ : std_logic;
signal \N__65282\ : std_logic;
signal \N__65281\ : std_logic;
signal \N__65280\ : std_logic;
signal \N__65273\ : std_logic;
signal \N__65272\ : std_logic;
signal \N__65271\ : std_logic;
signal \N__65264\ : std_logic;
signal \N__65263\ : std_logic;
signal \N__65262\ : std_logic;
signal \N__65255\ : std_logic;
signal \N__65254\ : std_logic;
signal \N__65253\ : std_logic;
signal \N__65246\ : std_logic;
signal \N__65245\ : std_logic;
signal \N__65244\ : std_logic;
signal \N__65237\ : std_logic;
signal \N__65236\ : std_logic;
signal \N__65235\ : std_logic;
signal \N__65228\ : std_logic;
signal \N__65227\ : std_logic;
signal \N__65226\ : std_logic;
signal \N__65219\ : std_logic;
signal \N__65218\ : std_logic;
signal \N__65217\ : std_logic;
signal \N__65210\ : std_logic;
signal \N__65209\ : std_logic;
signal \N__65208\ : std_logic;
signal \N__65201\ : std_logic;
signal \N__65200\ : std_logic;
signal \N__65199\ : std_logic;
signal \N__65192\ : std_logic;
signal \N__65191\ : std_logic;
signal \N__65190\ : std_logic;
signal \N__65183\ : std_logic;
signal \N__65182\ : std_logic;
signal \N__65181\ : std_logic;
signal \N__65174\ : std_logic;
signal \N__65173\ : std_logic;
signal \N__65172\ : std_logic;
signal \N__65165\ : std_logic;
signal \N__65164\ : std_logic;
signal \N__65163\ : std_logic;
signal \N__65156\ : std_logic;
signal \N__65155\ : std_logic;
signal \N__65154\ : std_logic;
signal \N__65147\ : std_logic;
signal \N__65146\ : std_logic;
signal \N__65145\ : std_logic;
signal \N__65138\ : std_logic;
signal \N__65137\ : std_logic;
signal \N__65136\ : std_logic;
signal \N__65129\ : std_logic;
signal \N__65128\ : std_logic;
signal \N__65127\ : std_logic;
signal \N__65120\ : std_logic;
signal \N__65119\ : std_logic;
signal \N__65118\ : std_logic;
signal \N__65111\ : std_logic;
signal \N__65110\ : std_logic;
signal \N__65109\ : std_logic;
signal \N__65102\ : std_logic;
signal \N__65101\ : std_logic;
signal \N__65100\ : std_logic;
signal \N__65093\ : std_logic;
signal \N__65092\ : std_logic;
signal \N__65091\ : std_logic;
signal \N__65084\ : std_logic;
signal \N__65083\ : std_logic;
signal \N__65082\ : std_logic;
signal \N__65075\ : std_logic;
signal \N__65074\ : std_logic;
signal \N__65073\ : std_logic;
signal \N__65066\ : std_logic;
signal \N__65065\ : std_logic;
signal \N__65064\ : std_logic;
signal \N__65057\ : std_logic;
signal \N__65056\ : std_logic;
signal \N__65055\ : std_logic;
signal \N__65048\ : std_logic;
signal \N__65047\ : std_logic;
signal \N__65046\ : std_logic;
signal \N__65039\ : std_logic;
signal \N__65038\ : std_logic;
signal \N__65037\ : std_logic;
signal \N__65030\ : std_logic;
signal \N__65029\ : std_logic;
signal \N__65028\ : std_logic;
signal \N__65021\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65019\ : std_logic;
signal \N__65012\ : std_logic;
signal \N__65011\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65003\ : std_logic;
signal \N__65002\ : std_logic;
signal \N__65001\ : std_logic;
signal \N__64984\ : std_logic;
signal \N__64981\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64977\ : std_logic;
signal \N__64974\ : std_logic;
signal \N__64971\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64963\ : std_logic;
signal \N__64962\ : std_logic;
signal \N__64959\ : std_logic;
signal \N__64956\ : std_logic;
signal \N__64951\ : std_logic;
signal \N__64948\ : std_logic;
signal \N__64947\ : std_logic;
signal \N__64944\ : std_logic;
signal \N__64941\ : std_logic;
signal \N__64936\ : std_logic;
signal \N__64933\ : std_logic;
signal \N__64932\ : std_logic;
signal \N__64929\ : std_logic;
signal \N__64926\ : std_logic;
signal \N__64921\ : std_logic;
signal \N__64918\ : std_logic;
signal \N__64917\ : std_logic;
signal \N__64914\ : std_logic;
signal \N__64911\ : std_logic;
signal \N__64906\ : std_logic;
signal \N__64903\ : std_logic;
signal \N__64902\ : std_logic;
signal \N__64899\ : std_logic;
signal \N__64896\ : std_logic;
signal \N__64891\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64887\ : std_logic;
signal \N__64884\ : std_logic;
signal \N__64881\ : std_logic;
signal \N__64876\ : std_logic;
signal \N__64873\ : std_logic;
signal \N__64870\ : std_logic;
signal \N__64869\ : std_logic;
signal \N__64868\ : std_logic;
signal \N__64865\ : std_logic;
signal \N__64862\ : std_logic;
signal \N__64859\ : std_logic;
signal \N__64858\ : std_logic;
signal \N__64857\ : std_logic;
signal \N__64856\ : std_logic;
signal \N__64855\ : std_logic;
signal \N__64854\ : std_logic;
signal \N__64853\ : std_logic;
signal \N__64852\ : std_logic;
signal \N__64851\ : std_logic;
signal \N__64850\ : std_logic;
signal \N__64849\ : std_logic;
signal \N__64848\ : std_logic;
signal \N__64847\ : std_logic;
signal \N__64846\ : std_logic;
signal \N__64845\ : std_logic;
signal \N__64844\ : std_logic;
signal \N__64841\ : std_logic;
signal \N__64836\ : std_logic;
signal \N__64833\ : std_logic;
signal \N__64830\ : std_logic;
signal \N__64829\ : std_logic;
signal \N__64828\ : std_logic;
signal \N__64825\ : std_logic;
signal \N__64824\ : std_logic;
signal \N__64823\ : std_logic;
signal \N__64820\ : std_logic;
signal \N__64819\ : std_logic;
signal \N__64816\ : std_logic;
signal \N__64815\ : std_logic;
signal \N__64812\ : std_logic;
signal \N__64811\ : std_logic;
signal \N__64808\ : std_logic;
signal \N__64807\ : std_logic;
signal \N__64804\ : std_logic;
signal \N__64803\ : std_logic;
signal \N__64800\ : std_logic;
signal \N__64799\ : std_logic;
signal \N__64796\ : std_logic;
signal \N__64795\ : std_logic;
signal \N__64792\ : std_logic;
signal \N__64789\ : std_logic;
signal \N__64788\ : std_logic;
signal \N__64785\ : std_logic;
signal \N__64784\ : std_logic;
signal \N__64781\ : std_logic;
signal \N__64780\ : std_logic;
signal \N__64777\ : std_logic;
signal \N__64774\ : std_logic;
signal \N__64767\ : std_logic;
signal \N__64764\ : std_logic;
signal \N__64761\ : std_logic;
signal \N__64758\ : std_logic;
signal \N__64755\ : std_logic;
signal \N__64752\ : std_logic;
signal \N__64749\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64733\ : std_logic;
signal \N__64732\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64730\ : std_logic;
signal \N__64729\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64727\ : std_logic;
signal \N__64712\ : std_logic;
signal \N__64697\ : std_logic;
signal \N__64696\ : std_logic;
signal \N__64695\ : std_logic;
signal \N__64694\ : std_logic;
signal \N__64693\ : std_logic;
signal \N__64684\ : std_logic;
signal \N__64677\ : std_logic;
signal \N__64676\ : std_logic;
signal \N__64673\ : std_logic;
signal \N__64670\ : std_logic;
signal \N__64667\ : std_logic;
signal \N__64666\ : std_logic;
signal \N__64663\ : std_logic;
signal \N__64660\ : std_logic;
signal \N__64657\ : std_logic;
signal \N__64654\ : std_logic;
signal \N__64651\ : std_logic;
signal \N__64648\ : std_logic;
signal \N__64645\ : std_logic;
signal \N__64642\ : std_logic;
signal \N__64641\ : std_logic;
signal \N__64638\ : std_logic;
signal \N__64637\ : std_logic;
signal \N__64634\ : std_logic;
signal \N__64633\ : std_logic;
signal \N__64630\ : std_logic;
signal \N__64629\ : std_logic;
signal \N__64626\ : std_logic;
signal \N__64621\ : std_logic;
signal \N__64618\ : std_logic;
signal \N__64617\ : std_logic;
signal \N__64616\ : std_logic;
signal \N__64613\ : std_logic;
signal \N__64610\ : std_logic;
signal \N__64601\ : std_logic;
signal \N__64592\ : std_logic;
signal \N__64587\ : std_logic;
signal \N__64570\ : std_logic;
signal \N__64567\ : std_logic;
signal \N__64564\ : std_logic;
signal \N__64561\ : std_logic;
signal \N__64558\ : std_logic;
signal \N__64557\ : std_logic;
signal \N__64554\ : std_logic;
signal \N__64551\ : std_logic;
signal \N__64542\ : std_logic;
signal \N__64537\ : std_logic;
signal \N__64534\ : std_logic;
signal \N__64531\ : std_logic;
signal \N__64528\ : std_logic;
signal \N__64521\ : std_logic;
signal \N__64518\ : std_logic;
signal \N__64513\ : std_logic;
signal \N__64510\ : std_logic;
signal \N__64501\ : std_logic;
signal \N__64498\ : std_logic;
signal \N__64497\ : std_logic;
signal \N__64494\ : std_logic;
signal \N__64491\ : std_logic;
signal \N__64488\ : std_logic;
signal \N__64483\ : std_logic;
signal \N__64480\ : std_logic;
signal \N__64479\ : std_logic;
signal \N__64476\ : std_logic;
signal \N__64473\ : std_logic;
signal \N__64470\ : std_logic;
signal \N__64467\ : std_logic;
signal \N__64462\ : std_logic;
signal \N__64459\ : std_logic;
signal \N__64458\ : std_logic;
signal \N__64457\ : std_logic;
signal \N__64454\ : std_logic;
signal \N__64451\ : std_logic;
signal \N__64448\ : std_logic;
signal \N__64447\ : std_logic;
signal \N__64444\ : std_logic;
signal \N__64441\ : std_logic;
signal \N__64438\ : std_logic;
signal \N__64435\ : std_logic;
signal \N__64432\ : std_logic;
signal \N__64427\ : std_logic;
signal \N__64424\ : std_logic;
signal \N__64417\ : std_logic;
signal \N__64416\ : std_logic;
signal \N__64413\ : std_logic;
signal \N__64410\ : std_logic;
signal \N__64407\ : std_logic;
signal \N__64404\ : std_logic;
signal \N__64401\ : std_logic;
signal \N__64398\ : std_logic;
signal \N__64393\ : std_logic;
signal \N__64392\ : std_logic;
signal \N__64389\ : std_logic;
signal \N__64386\ : std_logic;
signal \N__64381\ : std_logic;
signal \N__64378\ : std_logic;
signal \N__64377\ : std_logic;
signal \N__64374\ : std_logic;
signal \N__64371\ : std_logic;
signal \N__64366\ : std_logic;
signal \N__64363\ : std_logic;
signal \N__64360\ : std_logic;
signal \N__64359\ : std_logic;
signal \N__64356\ : std_logic;
signal \N__64353\ : std_logic;
signal \N__64348\ : std_logic;
signal \N__64345\ : std_logic;
signal \N__64342\ : std_logic;
signal \N__64341\ : std_logic;
signal \N__64338\ : std_logic;
signal \N__64335\ : std_logic;
signal \N__64330\ : std_logic;
signal \N__64327\ : std_logic;
signal \N__64326\ : std_logic;
signal \N__64323\ : std_logic;
signal \N__64320\ : std_logic;
signal \N__64317\ : std_logic;
signal \N__64314\ : std_logic;
signal \N__64311\ : std_logic;
signal \N__64306\ : std_logic;
signal \N__64303\ : std_logic;
signal \N__64302\ : std_logic;
signal \N__64299\ : std_logic;
signal \N__64296\ : std_logic;
signal \N__64291\ : std_logic;
signal \N__64288\ : std_logic;
signal \N__64285\ : std_logic;
signal \N__64284\ : std_logic;
signal \N__64281\ : std_logic;
signal \N__64278\ : std_logic;
signal \N__64273\ : std_logic;
signal \N__64270\ : std_logic;
signal \N__64269\ : std_logic;
signal \N__64266\ : std_logic;
signal \N__64263\ : std_logic;
signal \N__64260\ : std_logic;
signal \N__64255\ : std_logic;
signal \N__64252\ : std_logic;
signal \N__64249\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64243\ : std_logic;
signal \N__64240\ : std_logic;
signal \N__64237\ : std_logic;
signal \N__64234\ : std_logic;
signal \N__64231\ : std_logic;
signal \N__64228\ : std_logic;
signal \N__64227\ : std_logic;
signal \N__64224\ : std_logic;
signal \N__64221\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64219\ : std_logic;
signal \N__64218\ : std_logic;
signal \N__64217\ : std_logic;
signal \N__64216\ : std_logic;
signal \N__64211\ : std_logic;
signal \N__64206\ : std_logic;
signal \N__64203\ : std_logic;
signal \N__64198\ : std_logic;
signal \N__64189\ : std_logic;
signal \N__64186\ : std_logic;
signal \N__64183\ : std_logic;
signal \N__64180\ : std_logic;
signal \N__64179\ : std_logic;
signal \N__64176\ : std_logic;
signal \N__64173\ : std_logic;
signal \N__64168\ : std_logic;
signal \N__64167\ : std_logic;
signal \N__64164\ : std_logic;
signal \N__64163\ : std_logic;
signal \N__64162\ : std_logic;
signal \N__64161\ : std_logic;
signal \N__64154\ : std_logic;
signal \N__64151\ : std_logic;
signal \N__64148\ : std_logic;
signal \N__64143\ : std_logic;
signal \N__64138\ : std_logic;
signal \N__64135\ : std_logic;
signal \N__64132\ : std_logic;
signal \N__64129\ : std_logic;
signal \N__64126\ : std_logic;
signal \N__64123\ : std_logic;
signal \N__64120\ : std_logic;
signal \N__64117\ : std_logic;
signal \N__64114\ : std_logic;
signal \N__64111\ : std_logic;
signal \N__64110\ : std_logic;
signal \N__64109\ : std_logic;
signal \N__64102\ : std_logic;
signal \N__64101\ : std_logic;
signal \N__64098\ : std_logic;
signal \N__64097\ : std_logic;
signal \N__64096\ : std_logic;
signal \N__64095\ : std_logic;
signal \N__64092\ : std_logic;
signal \N__64091\ : std_logic;
signal \N__64090\ : std_logic;
signal \N__64089\ : std_logic;
signal \N__64088\ : std_logic;
signal \N__64085\ : std_logic;
signal \N__64080\ : std_logic;
signal \N__64079\ : std_logic;
signal \N__64078\ : std_logic;
signal \N__64077\ : std_logic;
signal \N__64076\ : std_logic;
signal \N__64067\ : std_logic;
signal \N__64066\ : std_logic;
signal \N__64065\ : std_logic;
signal \N__64062\ : std_logic;
signal \N__64059\ : std_logic;
signal \N__64054\ : std_logic;
signal \N__64051\ : std_logic;
signal \N__64050\ : std_logic;
signal \N__64049\ : std_logic;
signal \N__64048\ : std_logic;
signal \N__64041\ : std_logic;
signal \N__64038\ : std_logic;
signal \N__64035\ : std_logic;
signal \N__64034\ : std_logic;
signal \N__64033\ : std_logic;
signal \N__64032\ : std_logic;
signal \N__64031\ : std_logic;
signal \N__64030\ : std_logic;
signal \N__64029\ : std_logic;
signal \N__64026\ : std_logic;
signal \N__64025\ : std_logic;
signal \N__64024\ : std_logic;
signal \N__64023\ : std_logic;
signal \N__64022\ : std_logic;
signal \N__64017\ : std_logic;
signal \N__64012\ : std_logic;
signal \N__64011\ : std_logic;
signal \N__64008\ : std_logic;
signal \N__64007\ : std_logic;
signal \N__64006\ : std_logic;
signal \N__64001\ : std_logic;
signal \N__63998\ : std_logic;
signal \N__63995\ : std_logic;
signal \N__63994\ : std_logic;
signal \N__63993\ : std_logic;
signal \N__63992\ : std_logic;
signal \N__63991\ : std_logic;
signal \N__63990\ : std_logic;
signal \N__63989\ : std_logic;
signal \N__63988\ : std_logic;
signal \N__63987\ : std_logic;
signal \N__63986\ : std_logic;
signal \N__63985\ : std_logic;
signal \N__63980\ : std_logic;
signal \N__63973\ : std_logic;
signal \N__63970\ : std_logic;
signal \N__63967\ : std_logic;
signal \N__63966\ : std_logic;
signal \N__63963\ : std_logic;
signal \N__63960\ : std_logic;
signal \N__63959\ : std_logic;
signal \N__63956\ : std_logic;
signal \N__63951\ : std_logic;
signal \N__63946\ : std_logic;
signal \N__63941\ : std_logic;
signal \N__63936\ : std_logic;
signal \N__63931\ : std_logic;
signal \N__63928\ : std_logic;
signal \N__63923\ : std_logic;
signal \N__63920\ : std_logic;
signal \N__63911\ : std_logic;
signal \N__63910\ : std_logic;
signal \N__63909\ : std_logic;
signal \N__63908\ : std_logic;
signal \N__63905\ : std_logic;
signal \N__63902\ : std_logic;
signal \N__63899\ : std_logic;
signal \N__63896\ : std_logic;
signal \N__63893\ : std_logic;
signal \N__63890\ : std_logic;
signal \N__63889\ : std_logic;
signal \N__63888\ : std_logic;
signal \N__63885\ : std_logic;
signal \N__63882\ : std_logic;
signal \N__63879\ : std_logic;
signal \N__63876\ : std_logic;
signal \N__63873\ : std_logic;
signal \N__63868\ : std_logic;
signal \N__63865\ : std_logic;
signal \N__63860\ : std_logic;
signal \N__63853\ : std_logic;
signal \N__63848\ : std_logic;
signal \N__63845\ : std_logic;
signal \N__63836\ : std_logic;
signal \N__63827\ : std_logic;
signal \N__63822\ : std_logic;
signal \N__63815\ : std_logic;
signal \N__63802\ : std_logic;
signal \N__63799\ : std_logic;
signal \N__63784\ : std_logic;
signal \N__63783\ : std_logic;
signal \N__63782\ : std_logic;
signal \N__63781\ : std_logic;
signal \N__63780\ : std_logic;
signal \N__63779\ : std_logic;
signal \N__63778\ : std_logic;
signal \N__63777\ : std_logic;
signal \N__63774\ : std_logic;
signal \N__63771\ : std_logic;
signal \N__63770\ : std_logic;
signal \N__63769\ : std_logic;
signal \N__63768\ : std_logic;
signal \N__63767\ : std_logic;
signal \N__63766\ : std_logic;
signal \N__63765\ : std_logic;
signal \N__63764\ : std_logic;
signal \N__63763\ : std_logic;
signal \N__63762\ : std_logic;
signal \N__63761\ : std_logic;
signal \N__63760\ : std_logic;
signal \N__63757\ : std_logic;
signal \N__63756\ : std_logic;
signal \N__63753\ : std_logic;
signal \N__63752\ : std_logic;
signal \N__63749\ : std_logic;
signal \N__63748\ : std_logic;
signal \N__63745\ : std_logic;
signal \N__63744\ : std_logic;
signal \N__63743\ : std_logic;
signal \N__63742\ : std_logic;
signal \N__63741\ : std_logic;
signal \N__63740\ : std_logic;
signal \N__63739\ : std_logic;
signal \N__63738\ : std_logic;
signal \N__63737\ : std_logic;
signal \N__63736\ : std_logic;
signal \N__63735\ : std_logic;
signal \N__63732\ : std_logic;
signal \N__63727\ : std_logic;
signal \N__63726\ : std_logic;
signal \N__63725\ : std_logic;
signal \N__63724\ : std_logic;
signal \N__63723\ : std_logic;
signal \N__63722\ : std_logic;
signal \N__63719\ : std_logic;
signal \N__63718\ : std_logic;
signal \N__63717\ : std_logic;
signal \N__63714\ : std_logic;
signal \N__63711\ : std_logic;
signal \N__63708\ : std_logic;
signal \N__63705\ : std_logic;
signal \N__63702\ : std_logic;
signal \N__63699\ : std_logic;
signal \N__63696\ : std_logic;
signal \N__63693\ : std_logic;
signal \N__63690\ : std_logic;
signal \N__63687\ : std_logic;
signal \N__63670\ : std_logic;
signal \N__63667\ : std_logic;
signal \N__63656\ : std_logic;
signal \N__63655\ : std_logic;
signal \N__63654\ : std_logic;
signal \N__63651\ : std_logic;
signal \N__63650\ : std_logic;
signal \N__63649\ : std_logic;
signal \N__63648\ : std_logic;
signal \N__63645\ : std_logic;
signal \N__63644\ : std_logic;
signal \N__63643\ : std_logic;
signal \N__63642\ : std_logic;
signal \N__63637\ : std_logic;
signal \N__63634\ : std_logic;
signal \N__63631\ : std_logic;
signal \N__63628\ : std_logic;
signal \N__63625\ : std_logic;
signal \N__63622\ : std_logic;
signal \N__63619\ : std_logic;
signal \N__63618\ : std_logic;
signal \N__63617\ : std_logic;
signal \N__63614\ : std_logic;
signal \N__63613\ : std_logic;
signal \N__63612\ : std_logic;
signal \N__63611\ : std_logic;
signal \N__63610\ : std_logic;
signal \N__63609\ : std_logic;
signal \N__63608\ : std_logic;
signal \N__63607\ : std_logic;
signal \N__63606\ : std_logic;
signal \N__63605\ : std_logic;
signal \N__63604\ : std_logic;
signal \N__63603\ : std_logic;
signal \N__63602\ : std_logic;
signal \N__63601\ : std_logic;
signal \N__63598\ : std_logic;
signal \N__63597\ : std_logic;
signal \N__63596\ : std_logic;
signal \N__63595\ : std_logic;
signal \N__63594\ : std_logic;
signal \N__63589\ : std_logic;
signal \N__63580\ : std_logic;
signal \N__63571\ : std_logic;
signal \N__63568\ : std_logic;
signal \N__63559\ : std_logic;
signal \N__63554\ : std_logic;
signal \N__63551\ : std_logic;
signal \N__63548\ : std_logic;
signal \N__63545\ : std_logic;
signal \N__63542\ : std_logic;
signal \N__63541\ : std_logic;
signal \N__63540\ : std_logic;
signal \N__63539\ : std_logic;
signal \N__63536\ : std_logic;
signal \N__63529\ : std_logic;
signal \N__63528\ : std_logic;
signal \N__63527\ : std_logic;
signal \N__63526\ : std_logic;
signal \N__63525\ : std_logic;
signal \N__63514\ : std_logic;
signal \N__63511\ : std_logic;
signal \N__63506\ : std_logic;
signal \N__63505\ : std_logic;
signal \N__63504\ : std_logic;
signal \N__63501\ : std_logic;
signal \N__63498\ : std_logic;
signal \N__63495\ : std_logic;
signal \N__63494\ : std_logic;
signal \N__63493\ : std_logic;
signal \N__63492\ : std_logic;
signal \N__63491\ : std_logic;
signal \N__63490\ : std_logic;
signal \N__63489\ : std_logic;
signal \N__63488\ : std_logic;
signal \N__63487\ : std_logic;
signal \N__63486\ : std_logic;
signal \N__63485\ : std_logic;
signal \N__63484\ : std_logic;
signal \N__63483\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63479\ : std_logic;
signal \N__63474\ : std_logic;
signal \N__63469\ : std_logic;
signal \N__63466\ : std_logic;
signal \N__63457\ : std_logic;
signal \N__63454\ : std_logic;
signal \N__63451\ : std_logic;
signal \N__63448\ : std_logic;
signal \N__63445\ : std_logic;
signal \N__63438\ : std_logic;
signal \N__63421\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63415\ : std_logic;
signal \N__63412\ : std_logic;
signal \N__63407\ : std_logic;
signal \N__63402\ : std_logic;
signal \N__63397\ : std_logic;
signal \N__63394\ : std_logic;
signal \N__63393\ : std_logic;
signal \N__63390\ : std_logic;
signal \N__63383\ : std_logic;
signal \N__63382\ : std_logic;
signal \N__63381\ : std_logic;
signal \N__63380\ : std_logic;
signal \N__63379\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63373\ : std_logic;
signal \N__63366\ : std_logic;
signal \N__63359\ : std_logic;
signal \N__63358\ : std_logic;
signal \N__63357\ : std_logic;
signal \N__63354\ : std_logic;
signal \N__63349\ : std_logic;
signal \N__63346\ : std_logic;
signal \N__63341\ : std_logic;
signal \N__63338\ : std_logic;
signal \N__63331\ : std_logic;
signal \N__63320\ : std_logic;
signal \N__63317\ : std_logic;
signal \N__63314\ : std_logic;
signal \N__63305\ : std_logic;
signal \N__63300\ : std_logic;
signal \N__63291\ : std_logic;
signal \N__63288\ : std_logic;
signal \N__63285\ : std_logic;
signal \N__63282\ : std_logic;
signal \N__63279\ : std_logic;
signal \N__63270\ : std_logic;
signal \N__63267\ : std_logic;
signal \N__63260\ : std_logic;
signal \N__63255\ : std_logic;
signal \N__63240\ : std_logic;
signal \N__63229\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63205\ : std_logic;
signal \N__63204\ : std_logic;
signal \N__63201\ : std_logic;
signal \N__63200\ : std_logic;
signal \N__63197\ : std_logic;
signal \N__63196\ : std_logic;
signal \N__63195\ : std_logic;
signal \N__63194\ : std_logic;
signal \N__63191\ : std_logic;
signal \N__63190\ : std_logic;
signal \N__63189\ : std_logic;
signal \N__63188\ : std_logic;
signal \N__63185\ : std_logic;
signal \N__63182\ : std_logic;
signal \N__63177\ : std_logic;
signal \N__63174\ : std_logic;
signal \N__63173\ : std_logic;
signal \N__63170\ : std_logic;
signal \N__63167\ : std_logic;
signal \N__63164\ : std_logic;
signal \N__63163\ : std_logic;
signal \N__63162\ : std_logic;
signal \N__63157\ : std_logic;
signal \N__63152\ : std_logic;
signal \N__63149\ : std_logic;
signal \N__63146\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63140\ : std_logic;
signal \N__63133\ : std_logic;
signal \N__63128\ : std_logic;
signal \N__63125\ : std_logic;
signal \N__63122\ : std_logic;
signal \N__63119\ : std_logic;
signal \N__63114\ : std_logic;
signal \N__63111\ : std_logic;
signal \N__63110\ : std_logic;
signal \N__63105\ : std_logic;
signal \N__63100\ : std_logic;
signal \N__63097\ : std_logic;
signal \N__63094\ : std_logic;
signal \N__63085\ : std_logic;
signal \N__63084\ : std_logic;
signal \N__63083\ : std_logic;
signal \N__63082\ : std_logic;
signal \N__63081\ : std_logic;
signal \N__63080\ : std_logic;
signal \N__63079\ : std_logic;
signal \N__63078\ : std_logic;
signal \N__63077\ : std_logic;
signal \N__63076\ : std_logic;
signal \N__63075\ : std_logic;
signal \N__63074\ : std_logic;
signal \N__63073\ : std_logic;
signal \N__63072\ : std_logic;
signal \N__63071\ : std_logic;
signal \N__63070\ : std_logic;
signal \N__63067\ : std_logic;
signal \N__63066\ : std_logic;
signal \N__63061\ : std_logic;
signal \N__63060\ : std_logic;
signal \N__63059\ : std_logic;
signal \N__63058\ : std_logic;
signal \N__63057\ : std_logic;
signal \N__63056\ : std_logic;
signal \N__63055\ : std_logic;
signal \N__63052\ : std_logic;
signal \N__63051\ : std_logic;
signal \N__63050\ : std_logic;
signal \N__63049\ : std_logic;
signal \N__63048\ : std_logic;
signal \N__63047\ : std_logic;
signal \N__63046\ : std_logic;
signal \N__63045\ : std_logic;
signal \N__63042\ : std_logic;
signal \N__63039\ : std_logic;
signal \N__63034\ : std_logic;
signal \N__63031\ : std_logic;
signal \N__63030\ : std_logic;
signal \N__63029\ : std_logic;
signal \N__63028\ : std_logic;
signal \N__63027\ : std_logic;
signal \N__63024\ : std_logic;
signal \N__63021\ : std_logic;
signal \N__63018\ : std_logic;
signal \N__63015\ : std_logic;
signal \N__63012\ : std_logic;
signal \N__63003\ : std_logic;
signal \N__63000\ : std_logic;
signal \N__62991\ : std_logic;
signal \N__62986\ : std_logic;
signal \N__62983\ : std_logic;
signal \N__62980\ : std_logic;
signal \N__62973\ : std_logic;
signal \N__62970\ : std_logic;
signal \N__62969\ : std_logic;
signal \N__62964\ : std_logic;
signal \N__62957\ : std_logic;
signal \N__62954\ : std_logic;
signal \N__62949\ : std_logic;
signal \N__62944\ : std_logic;
signal \N__62943\ : std_logic;
signal \N__62940\ : std_logic;
signal \N__62937\ : std_logic;
signal \N__62936\ : std_logic;
signal \N__62935\ : std_logic;
signal \N__62934\ : std_logic;
signal \N__62933\ : std_logic;
signal \N__62932\ : std_logic;
signal \N__62931\ : std_logic;
signal \N__62930\ : std_logic;
signal \N__62927\ : std_logic;
signal \N__62924\ : std_logic;
signal \N__62913\ : std_logic;
signal \N__62908\ : std_logic;
signal \N__62907\ : std_logic;
signal \N__62906\ : std_logic;
signal \N__62905\ : std_logic;
signal \N__62902\ : std_logic;
signal \N__62899\ : std_logic;
signal \N__62896\ : std_logic;
signal \N__62891\ : std_logic;
signal \N__62884\ : std_logic;
signal \N__62881\ : std_logic;
signal \N__62878\ : std_logic;
signal \N__62875\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62863\ : std_logic;
signal \N__62858\ : std_logic;
signal \N__62849\ : std_logic;
signal \N__62844\ : std_logic;
signal \N__62841\ : std_logic;
signal \N__62836\ : std_logic;
signal \N__62831\ : std_logic;
signal \N__62822\ : std_logic;
signal \N__62803\ : std_logic;
signal \N__62800\ : std_logic;
signal \N__62797\ : std_logic;
signal \N__62794\ : std_logic;
signal \N__62791\ : std_logic;
signal \N__62790\ : std_logic;
signal \N__62789\ : std_logic;
signal \N__62788\ : std_logic;
signal \N__62785\ : std_logic;
signal \N__62784\ : std_logic;
signal \N__62781\ : std_logic;
signal \N__62780\ : std_logic;
signal \N__62779\ : std_logic;
signal \N__62776\ : std_logic;
signal \N__62775\ : std_logic;
signal \N__62772\ : std_logic;
signal \N__62769\ : std_logic;
signal \N__62766\ : std_logic;
signal \N__62763\ : std_logic;
signal \N__62760\ : std_logic;
signal \N__62757\ : std_logic;
signal \N__62754\ : std_logic;
signal \N__62751\ : std_logic;
signal \N__62748\ : std_logic;
signal \N__62743\ : std_logic;
signal \N__62740\ : std_logic;
signal \N__62737\ : std_logic;
signal \N__62734\ : std_logic;
signal \N__62731\ : std_logic;
signal \N__62728\ : std_logic;
signal \N__62727\ : std_logic;
signal \N__62724\ : std_logic;
signal \N__62721\ : std_logic;
signal \N__62716\ : std_logic;
signal \N__62713\ : std_logic;
signal \N__62708\ : std_logic;
signal \N__62705\ : std_logic;
signal \N__62692\ : std_logic;
signal \N__62691\ : std_logic;
signal \N__62690\ : std_logic;
signal \N__62689\ : std_logic;
signal \N__62686\ : std_logic;
signal \N__62685\ : std_logic;
signal \N__62682\ : std_logic;
signal \N__62679\ : std_logic;
signal \N__62678\ : std_logic;
signal \N__62677\ : std_logic;
signal \N__62676\ : std_logic;
signal \N__62675\ : std_logic;
signal \N__62674\ : std_logic;
signal \N__62673\ : std_logic;
signal \N__62672\ : std_logic;
signal \N__62671\ : std_logic;
signal \N__62670\ : std_logic;
signal \N__62667\ : std_logic;
signal \N__62664\ : std_logic;
signal \N__62663\ : std_logic;
signal \N__62662\ : std_logic;
signal \N__62661\ : std_logic;
signal \N__62660\ : std_logic;
signal \N__62659\ : std_logic;
signal \N__62658\ : std_logic;
signal \N__62657\ : std_logic;
signal \N__62656\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62654\ : std_logic;
signal \N__62653\ : std_logic;
signal \N__62652\ : std_logic;
signal \N__62649\ : std_logic;
signal \N__62648\ : std_logic;
signal \N__62647\ : std_logic;
signal \N__62646\ : std_logic;
signal \N__62645\ : std_logic;
signal \N__62638\ : std_logic;
signal \N__62637\ : std_logic;
signal \N__62634\ : std_logic;
signal \N__62633\ : std_logic;
signal \N__62632\ : std_logic;
signal \N__62631\ : std_logic;
signal \N__62630\ : std_logic;
signal \N__62629\ : std_logic;
signal \N__62628\ : std_logic;
signal \N__62627\ : std_logic;
signal \N__62626\ : std_logic;
signal \N__62625\ : std_logic;
signal \N__62624\ : std_logic;
signal \N__62623\ : std_logic;
signal \N__62622\ : std_logic;
signal \N__62621\ : std_logic;
signal \N__62620\ : std_logic;
signal \N__62619\ : std_logic;
signal \N__62618\ : std_logic;
signal \N__62617\ : std_logic;
signal \N__62616\ : std_logic;
signal \N__62615\ : std_logic;
signal \N__62612\ : std_logic;
signal \N__62611\ : std_logic;
signal \N__62610\ : std_logic;
signal \N__62609\ : std_logic;
signal \N__62608\ : std_logic;
signal \N__62607\ : std_logic;
signal \N__62606\ : std_logic;
signal \N__62605\ : std_logic;
signal \N__62604\ : std_logic;
signal \N__62603\ : std_logic;
signal \N__62602\ : std_logic;
signal \N__62601\ : std_logic;
signal \N__62600\ : std_logic;
signal \N__62599\ : std_logic;
signal \N__62598\ : std_logic;
signal \N__62597\ : std_logic;
signal \N__62596\ : std_logic;
signal \N__62595\ : std_logic;
signal \N__62588\ : std_logic;
signal \N__62585\ : std_logic;
signal \N__62582\ : std_logic;
signal \N__62579\ : std_logic;
signal \N__62576\ : std_logic;
signal \N__62573\ : std_logic;
signal \N__62572\ : std_logic;
signal \N__62571\ : std_logic;
signal \N__62570\ : std_logic;
signal \N__62569\ : std_logic;
signal \N__62568\ : std_logic;
signal \N__62567\ : std_logic;
signal \N__62566\ : std_logic;
signal \N__62565\ : std_logic;
signal \N__62564\ : std_logic;
signal \N__62561\ : std_logic;
signal \N__62548\ : std_logic;
signal \N__62531\ : std_logic;
signal \N__62530\ : std_logic;
signal \N__62529\ : std_logic;
signal \N__62528\ : std_logic;
signal \N__62527\ : std_logic;
signal \N__62526\ : std_logic;
signal \N__62525\ : std_logic;
signal \N__62524\ : std_logic;
signal \N__62523\ : std_logic;
signal \N__62522\ : std_logic;
signal \N__62521\ : std_logic;
signal \N__62516\ : std_logic;
signal \N__62513\ : std_logic;
signal \N__62510\ : std_logic;
signal \N__62507\ : std_logic;
signal \N__62504\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62486\ : std_logic;
signal \N__62485\ : std_logic;
signal \N__62482\ : std_logic;
signal \N__62481\ : std_logic;
signal \N__62480\ : std_logic;
signal \N__62463\ : std_logic;
signal \N__62460\ : std_logic;
signal \N__62451\ : std_logic;
signal \N__62450\ : std_logic;
signal \N__62449\ : std_logic;
signal \N__62446\ : std_logic;
signal \N__62443\ : std_logic;
signal \N__62440\ : std_logic;
signal \N__62435\ : std_logic;
signal \N__62432\ : std_logic;
signal \N__62429\ : std_logic;
signal \N__62428\ : std_logic;
signal \N__62427\ : std_logic;
signal \N__62426\ : std_logic;
signal \N__62423\ : std_logic;
signal \N__62422\ : std_logic;
signal \N__62421\ : std_logic;
signal \N__62418\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62406\ : std_logic;
signal \N__62403\ : std_logic;
signal \N__62392\ : std_logic;
signal \N__62385\ : std_logic;
signal \N__62380\ : std_logic;
signal \N__62373\ : std_logic;
signal \N__62370\ : std_logic;
signal \N__62369\ : std_logic;
signal \N__62368\ : std_logic;
signal \N__62361\ : std_logic;
signal \N__62358\ : std_logic;
signal \N__62355\ : std_logic;
signal \N__62338\ : std_logic;
signal \N__62335\ : std_logic;
signal \N__62332\ : std_logic;
signal \N__62327\ : std_logic;
signal \N__62324\ : std_logic;
signal \N__62321\ : std_logic;
signal \N__62316\ : std_logic;
signal \N__62313\ : std_logic;
signal \N__62308\ : std_logic;
signal \N__62301\ : std_logic;
signal \N__62298\ : std_logic;
signal \N__62297\ : std_logic;
signal \N__62296\ : std_logic;
signal \N__62295\ : std_logic;
signal \N__62294\ : std_logic;
signal \N__62293\ : std_logic;
signal \N__62292\ : std_logic;
signal \N__62291\ : std_logic;
signal \N__62290\ : std_logic;
signal \N__62285\ : std_logic;
signal \N__62276\ : std_logic;
signal \N__62273\ : std_logic;
signal \N__62260\ : std_logic;
signal \N__62243\ : std_logic;
signal \N__62242\ : std_logic;
signal \N__62241\ : std_logic;
signal \N__62240\ : std_logic;
signal \N__62237\ : std_logic;
signal \N__62232\ : std_logic;
signal \N__62227\ : std_logic;
signal \N__62218\ : std_logic;
signal \N__62215\ : std_logic;
signal \N__62212\ : std_logic;
signal \N__62205\ : std_logic;
signal \N__62200\ : std_logic;
signal \N__62197\ : std_logic;
signal \N__62192\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62184\ : std_logic;
signal \N__62179\ : std_logic;
signal \N__62176\ : std_logic;
signal \N__62171\ : std_logic;
signal \N__62164\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62154\ : std_logic;
signal \N__62145\ : std_logic;
signal \N__62138\ : std_logic;
signal \N__62113\ : std_logic;
signal \N__62110\ : std_logic;
signal \N__62107\ : std_logic;
signal \N__62104\ : std_logic;
signal \N__62101\ : std_logic;
signal \N__62100\ : std_logic;
signal \N__62097\ : std_logic;
signal \N__62094\ : std_logic;
signal \N__62093\ : std_logic;
signal \N__62092\ : std_logic;
signal \N__62087\ : std_logic;
signal \N__62086\ : std_logic;
signal \N__62083\ : std_logic;
signal \N__62080\ : std_logic;
signal \N__62079\ : std_logic;
signal \N__62076\ : std_logic;
signal \N__62073\ : std_logic;
signal \N__62070\ : std_logic;
signal \N__62065\ : std_logic;
signal \N__62060\ : std_logic;
signal \N__62057\ : std_logic;
signal \N__62056\ : std_logic;
signal \N__62053\ : std_logic;
signal \N__62050\ : std_logic;
signal \N__62047\ : std_logic;
signal \N__62044\ : std_logic;
signal \N__62041\ : std_logic;
signal \N__62038\ : std_logic;
signal \N__62033\ : std_logic;
signal \N__62030\ : std_logic;
signal \N__62025\ : std_logic;
signal \N__62022\ : std_logic;
signal \N__62019\ : std_logic;
signal \N__62014\ : std_logic;
signal \N__62013\ : std_logic;
signal \N__62012\ : std_logic;
signal \N__62011\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62009\ : std_logic;
signal \N__62008\ : std_logic;
signal \N__62007\ : std_logic;
signal \N__62006\ : std_logic;
signal \N__62005\ : std_logic;
signal \N__62004\ : std_logic;
signal \N__62003\ : std_logic;
signal \N__62002\ : std_logic;
signal \N__62001\ : std_logic;
signal \N__62000\ : std_logic;
signal \N__61999\ : std_logic;
signal \N__61998\ : std_logic;
signal \N__61997\ : std_logic;
signal \N__61996\ : std_logic;
signal \N__61995\ : std_logic;
signal \N__61994\ : std_logic;
signal \N__61993\ : std_logic;
signal \N__61992\ : std_logic;
signal \N__61991\ : std_logic;
signal \N__61990\ : std_logic;
signal \N__61989\ : std_logic;
signal \N__61988\ : std_logic;
signal \N__61987\ : std_logic;
signal \N__61986\ : std_logic;
signal \N__61985\ : std_logic;
signal \N__61984\ : std_logic;
signal \N__61983\ : std_logic;
signal \N__61982\ : std_logic;
signal \N__61981\ : std_logic;
signal \N__61980\ : std_logic;
signal \N__61979\ : std_logic;
signal \N__61978\ : std_logic;
signal \N__61977\ : std_logic;
signal \N__61976\ : std_logic;
signal \N__61975\ : std_logic;
signal \N__61974\ : std_logic;
signal \N__61973\ : std_logic;
signal \N__61972\ : std_logic;
signal \N__61971\ : std_logic;
signal \N__61970\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61968\ : std_logic;
signal \N__61967\ : std_logic;
signal \N__61966\ : std_logic;
signal \N__61965\ : std_logic;
signal \N__61964\ : std_logic;
signal \N__61963\ : std_logic;
signal \N__61962\ : std_logic;
signal \N__61961\ : std_logic;
signal \N__61960\ : std_logic;
signal \N__61959\ : std_logic;
signal \N__61958\ : std_logic;
signal \N__61957\ : std_logic;
signal \N__61956\ : std_logic;
signal \N__61955\ : std_logic;
signal \N__61954\ : std_logic;
signal \N__61953\ : std_logic;
signal \N__61952\ : std_logic;
signal \N__61951\ : std_logic;
signal \N__61950\ : std_logic;
signal \N__61949\ : std_logic;
signal \N__61948\ : std_logic;
signal \N__61947\ : std_logic;
signal \N__61946\ : std_logic;
signal \N__61945\ : std_logic;
signal \N__61944\ : std_logic;
signal \N__61943\ : std_logic;
signal \N__61942\ : std_logic;
signal \N__61941\ : std_logic;
signal \N__61940\ : std_logic;
signal \N__61939\ : std_logic;
signal \N__61938\ : std_logic;
signal \N__61937\ : std_logic;
signal \N__61936\ : std_logic;
signal \N__61935\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61933\ : std_logic;
signal \N__61932\ : std_logic;
signal \N__61931\ : std_logic;
signal \N__61930\ : std_logic;
signal \N__61929\ : std_logic;
signal \N__61928\ : std_logic;
signal \N__61927\ : std_logic;
signal \N__61926\ : std_logic;
signal \N__61925\ : std_logic;
signal \N__61924\ : std_logic;
signal \N__61923\ : std_logic;
signal \N__61922\ : std_logic;
signal \N__61921\ : std_logic;
signal \N__61920\ : std_logic;
signal \N__61919\ : std_logic;
signal \N__61918\ : std_logic;
signal \N__61917\ : std_logic;
signal \N__61916\ : std_logic;
signal \N__61915\ : std_logic;
signal \N__61914\ : std_logic;
signal \N__61913\ : std_logic;
signal \N__61912\ : std_logic;
signal \N__61911\ : std_logic;
signal \N__61910\ : std_logic;
signal \N__61909\ : std_logic;
signal \N__61908\ : std_logic;
signal \N__61907\ : std_logic;
signal \N__61906\ : std_logic;
signal \N__61905\ : std_logic;
signal \N__61904\ : std_logic;
signal \N__61903\ : std_logic;
signal \N__61902\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61900\ : std_logic;
signal \N__61899\ : std_logic;
signal \N__61898\ : std_logic;
signal \N__61897\ : std_logic;
signal \N__61896\ : std_logic;
signal \N__61895\ : std_logic;
signal \N__61894\ : std_logic;
signal \N__61893\ : std_logic;
signal \N__61892\ : std_logic;
signal \N__61891\ : std_logic;
signal \N__61890\ : std_logic;
signal \N__61889\ : std_logic;
signal \N__61888\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61886\ : std_logic;
signal \N__61885\ : std_logic;
signal \N__61884\ : std_logic;
signal \N__61883\ : std_logic;
signal \N__61882\ : std_logic;
signal \N__61881\ : std_logic;
signal \N__61880\ : std_logic;
signal \N__61879\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61877\ : std_logic;
signal \N__61876\ : std_logic;
signal \N__61875\ : std_logic;
signal \N__61874\ : std_logic;
signal \N__61873\ : std_logic;
signal \N__61872\ : std_logic;
signal \N__61871\ : std_logic;
signal \N__61870\ : std_logic;
signal \N__61869\ : std_logic;
signal \N__61868\ : std_logic;
signal \N__61867\ : std_logic;
signal \N__61866\ : std_logic;
signal \N__61865\ : std_logic;
signal \N__61864\ : std_logic;
signal \N__61863\ : std_logic;
signal \N__61862\ : std_logic;
signal \N__61861\ : std_logic;
signal \N__61860\ : std_logic;
signal \N__61859\ : std_logic;
signal \N__61858\ : std_logic;
signal \N__61857\ : std_logic;
signal \N__61856\ : std_logic;
signal \N__61855\ : std_logic;
signal \N__61854\ : std_logic;
signal \N__61853\ : std_logic;
signal \N__61852\ : std_logic;
signal \N__61851\ : std_logic;
signal \N__61850\ : std_logic;
signal \N__61849\ : std_logic;
signal \N__61848\ : std_logic;
signal \N__61847\ : std_logic;
signal \N__61846\ : std_logic;
signal \N__61845\ : std_logic;
signal \N__61844\ : std_logic;
signal \N__61843\ : std_logic;
signal \N__61842\ : std_logic;
signal \N__61841\ : std_logic;
signal \N__61840\ : std_logic;
signal \N__61839\ : std_logic;
signal \N__61838\ : std_logic;
signal \N__61837\ : std_logic;
signal \N__61836\ : std_logic;
signal \N__61835\ : std_logic;
signal \N__61834\ : std_logic;
signal \N__61833\ : std_logic;
signal \N__61832\ : std_logic;
signal \N__61831\ : std_logic;
signal \N__61830\ : std_logic;
signal \N__61829\ : std_logic;
signal \N__61828\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61826\ : std_logic;
signal \N__61825\ : std_logic;
signal \N__61824\ : std_logic;
signal \N__61441\ : std_logic;
signal \N__61438\ : std_logic;
signal \N__61437\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61431\ : std_logic;
signal \N__61428\ : std_logic;
signal \N__61425\ : std_logic;
signal \N__61420\ : std_logic;
signal \N__61417\ : std_logic;
signal \N__61414\ : std_logic;
signal \N__61413\ : std_logic;
signal \N__61412\ : std_logic;
signal \N__61411\ : std_logic;
signal \N__61410\ : std_logic;
signal \N__61409\ : std_logic;
signal \N__61408\ : std_logic;
signal \N__61407\ : std_logic;
signal \N__61406\ : std_logic;
signal \N__61405\ : std_logic;
signal \N__61402\ : std_logic;
signal \N__61401\ : std_logic;
signal \N__61400\ : std_logic;
signal \N__61399\ : std_logic;
signal \N__61398\ : std_logic;
signal \N__61397\ : std_logic;
signal \N__61396\ : std_logic;
signal \N__61395\ : std_logic;
signal \N__61394\ : std_logic;
signal \N__61391\ : std_logic;
signal \N__61390\ : std_logic;
signal \N__61387\ : std_logic;
signal \N__61384\ : std_logic;
signal \N__61383\ : std_logic;
signal \N__61382\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61380\ : std_logic;
signal \N__61379\ : std_logic;
signal \N__61376\ : std_logic;
signal \N__61375\ : std_logic;
signal \N__61374\ : std_logic;
signal \N__61373\ : std_logic;
signal \N__61370\ : std_logic;
signal \N__61367\ : std_logic;
signal \N__61364\ : std_logic;
signal \N__61363\ : std_logic;
signal \N__61362\ : std_logic;
signal \N__61359\ : std_logic;
signal \N__61356\ : std_logic;
signal \N__61353\ : std_logic;
signal \N__61352\ : std_logic;
signal \N__61349\ : std_logic;
signal \N__61348\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61344\ : std_logic;
signal \N__61339\ : std_logic;
signal \N__61336\ : std_logic;
signal \N__61333\ : std_logic;
signal \N__61330\ : std_logic;
signal \N__61327\ : std_logic;
signal \N__61322\ : std_logic;
signal \N__61319\ : std_logic;
signal \N__61316\ : std_logic;
signal \N__61313\ : std_logic;
signal \N__61310\ : std_logic;
signal \N__61307\ : std_logic;
signal \N__61304\ : std_logic;
signal \N__61301\ : std_logic;
signal \N__61300\ : std_logic;
signal \N__61297\ : std_logic;
signal \N__61292\ : std_logic;
signal \N__61291\ : std_logic;
signal \N__61288\ : std_logic;
signal \N__61281\ : std_logic;
signal \N__61276\ : std_logic;
signal \N__61269\ : std_logic;
signal \N__61268\ : std_logic;
signal \N__61267\ : std_logic;
signal \N__61264\ : std_logic;
signal \N__61261\ : std_logic;
signal \N__61260\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61254\ : std_logic;
signal \N__61253\ : std_logic;
signal \N__61248\ : std_logic;
signal \N__61245\ : std_logic;
signal \N__61242\ : std_logic;
signal \N__61233\ : std_logic;
signal \N__61232\ : std_logic;
signal \N__61231\ : std_logic;
signal \N__61226\ : std_logic;
signal \N__61223\ : std_logic;
signal \N__61218\ : std_logic;
signal \N__61215\ : std_logic;
signal \N__61212\ : std_logic;
signal \N__61207\ : std_logic;
signal \N__61204\ : std_logic;
signal \N__61201\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61189\ : std_logic;
signal \N__61184\ : std_logic;
signal \N__61183\ : std_logic;
signal \N__61182\ : std_logic;
signal \N__61179\ : std_logic;
signal \N__61178\ : std_logic;
signal \N__61175\ : std_logic;
signal \N__61172\ : std_logic;
signal \N__61169\ : std_logic;
signal \N__61160\ : std_logic;
signal \N__61157\ : std_logic;
signal \N__61154\ : std_logic;
signal \N__61141\ : std_logic;
signal \N__61130\ : std_logic;
signal \N__61121\ : std_logic;
signal \N__61102\ : std_logic;
signal \N__61099\ : std_logic;
signal \N__61096\ : std_logic;
signal \N__61095\ : std_logic;
signal \N__61092\ : std_logic;
signal \N__61089\ : std_logic;
signal \N__61086\ : std_logic;
signal \N__61083\ : std_logic;
signal \N__61080\ : std_logic;
signal \N__61075\ : std_logic;
signal \N__61072\ : std_logic;
signal \N__61069\ : std_logic;
signal \N__61066\ : std_logic;
signal \N__61063\ : std_logic;
signal \N__61060\ : std_logic;
signal \N__61057\ : std_logic;
signal \N__61056\ : std_logic;
signal \N__61055\ : std_logic;
signal \N__61054\ : std_logic;
signal \N__61053\ : std_logic;
signal \N__61052\ : std_logic;
signal \N__61051\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61042\ : std_logic;
signal \N__61037\ : std_logic;
signal \N__61036\ : std_logic;
signal \N__61035\ : std_logic;
signal \N__61034\ : std_logic;
signal \N__61033\ : std_logic;
signal \N__61032\ : std_logic;
signal \N__61029\ : std_logic;
signal \N__61026\ : std_logic;
signal \N__61025\ : std_logic;
signal \N__61024\ : std_logic;
signal \N__61023\ : std_logic;
signal \N__61022\ : std_logic;
signal \N__61021\ : std_logic;
signal \N__61020\ : std_logic;
signal \N__61019\ : std_logic;
signal \N__61018\ : std_logic;
signal \N__61017\ : std_logic;
signal \N__61014\ : std_logic;
signal \N__61013\ : std_logic;
signal \N__61010\ : std_logic;
signal \N__61007\ : std_logic;
signal \N__61004\ : std_logic;
signal \N__60995\ : std_logic;
signal \N__60994\ : std_logic;
signal \N__60993\ : std_logic;
signal \N__60992\ : std_logic;
signal \N__60991\ : std_logic;
signal \N__60990\ : std_logic;
signal \N__60989\ : std_logic;
signal \N__60986\ : std_logic;
signal \N__60981\ : std_logic;
signal \N__60980\ : std_logic;
signal \N__60979\ : std_logic;
signal \N__60978\ : std_logic;
signal \N__60977\ : std_logic;
signal \N__60976\ : std_logic;
signal \N__60975\ : std_logic;
signal \N__60970\ : std_logic;
signal \N__60963\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60957\ : std_logic;
signal \N__60956\ : std_logic;
signal \N__60955\ : std_logic;
signal \N__60954\ : std_logic;
signal \N__60953\ : std_logic;
signal \N__60952\ : std_logic;
signal \N__60949\ : std_logic;
signal \N__60948\ : std_logic;
signal \N__60945\ : std_logic;
signal \N__60942\ : std_logic;
signal \N__60939\ : std_logic;
signal \N__60932\ : std_logic;
signal \N__60929\ : std_logic;
signal \N__60926\ : std_logic;
signal \N__60921\ : std_logic;
signal \N__60918\ : std_logic;
signal \N__60915\ : std_logic;
signal \N__60912\ : std_logic;
signal \N__60909\ : std_logic;
signal \N__60906\ : std_logic;
signal \N__60903\ : std_logic;
signal \N__60902\ : std_logic;
signal \N__60899\ : std_logic;
signal \N__60894\ : std_logic;
signal \N__60889\ : std_logic;
signal \N__60884\ : std_logic;
signal \N__60881\ : std_logic;
signal \N__60880\ : std_logic;
signal \N__60879\ : std_logic;
signal \N__60876\ : std_logic;
signal \N__60871\ : std_logic;
signal \N__60866\ : std_logic;
signal \N__60865\ : std_logic;
signal \N__60862\ : std_logic;
signal \N__60859\ : std_logic;
signal \N__60856\ : std_logic;
signal \N__60853\ : std_logic;
signal \N__60850\ : std_logic;
signal \N__60847\ : std_logic;
signal \N__60842\ : std_logic;
signal \N__60837\ : std_logic;
signal \N__60834\ : std_logic;
signal \N__60831\ : std_logic;
signal \N__60822\ : std_logic;
signal \N__60819\ : std_logic;
signal \N__60810\ : std_logic;
signal \N__60807\ : std_logic;
signal \N__60804\ : std_logic;
signal \N__60801\ : std_logic;
signal \N__60794\ : std_logic;
signal \N__60793\ : std_logic;
signal \N__60792\ : std_logic;
signal \N__60789\ : std_logic;
signal \N__60786\ : std_logic;
signal \N__60781\ : std_logic;
signal \N__60778\ : std_logic;
signal \N__60775\ : std_logic;
signal \N__60770\ : std_logic;
signal \N__60757\ : std_logic;
signal \N__60750\ : std_logic;
signal \N__60747\ : std_logic;
signal \N__60742\ : std_logic;
signal \N__60721\ : std_logic;
signal \N__60718\ : std_logic;
signal \N__60715\ : std_logic;
signal \N__60712\ : std_logic;
signal \N__60709\ : std_logic;
signal \N__60706\ : std_logic;
signal \N__60703\ : std_logic;
signal \N__60700\ : std_logic;
signal \N__60697\ : std_logic;
signal \N__60694\ : std_logic;
signal \N__60691\ : std_logic;
signal \N__60690\ : std_logic;
signal \N__60689\ : std_logic;
signal \N__60686\ : std_logic;
signal \N__60681\ : std_logic;
signal \N__60676\ : std_logic;
signal \N__60673\ : std_logic;
signal \N__60670\ : std_logic;
signal \N__60669\ : std_logic;
signal \N__60668\ : std_logic;
signal \N__60667\ : std_logic;
signal \N__60666\ : std_logic;
signal \N__60665\ : std_logic;
signal \N__60664\ : std_logic;
signal \N__60663\ : std_logic;
signal \N__60660\ : std_logic;
signal \N__60657\ : std_logic;
signal \N__60650\ : std_logic;
signal \N__60649\ : std_logic;
signal \N__60648\ : std_logic;
signal \N__60647\ : std_logic;
signal \N__60646\ : std_logic;
signal \N__60643\ : std_logic;
signal \N__60642\ : std_logic;
signal \N__60641\ : std_logic;
signal \N__60640\ : std_logic;
signal \N__60637\ : std_logic;
signal \N__60636\ : std_logic;
signal \N__60635\ : std_logic;
signal \N__60632\ : std_logic;
signal \N__60631\ : std_logic;
signal \N__60628\ : std_logic;
signal \N__60627\ : std_logic;
signal \N__60624\ : std_logic;
signal \N__60621\ : std_logic;
signal \N__60620\ : std_logic;
signal \N__60619\ : std_logic;
signal \N__60616\ : std_logic;
signal \N__60615\ : std_logic;
signal \N__60612\ : std_logic;
signal \N__60611\ : std_logic;
signal \N__60610\ : std_logic;
signal \N__60609\ : std_logic;
signal \N__60604\ : std_logic;
signal \N__60603\ : std_logic;
signal \N__60602\ : std_logic;
signal \N__60601\ : std_logic;
signal \N__60600\ : std_logic;
signal \N__60599\ : std_logic;
signal \N__60598\ : std_logic;
signal \N__60597\ : std_logic;
signal \N__60596\ : std_logic;
signal \N__60595\ : std_logic;
signal \N__60594\ : std_logic;
signal \N__60593\ : std_logic;
signal \N__60592\ : std_logic;
signal \N__60591\ : std_logic;
signal \N__60590\ : std_logic;
signal \N__60589\ : std_logic;
signal \N__60588\ : std_logic;
signal \N__60587\ : std_logic;
signal \N__60584\ : std_logic;
signal \N__60579\ : std_logic;
signal \N__60576\ : std_logic;
signal \N__60573\ : std_logic;
signal \N__60568\ : std_logic;
signal \N__60565\ : std_logic;
signal \N__60564\ : std_logic;
signal \N__60561\ : std_logic;
signal \N__60558\ : std_logic;
signal \N__60555\ : std_logic;
signal \N__60550\ : std_logic;
signal \N__60547\ : std_logic;
signal \N__60546\ : std_logic;
signal \N__60545\ : std_logic;
signal \N__60544\ : std_logic;
signal \N__60543\ : std_logic;
signal \N__60540\ : std_logic;
signal \N__60537\ : std_logic;
signal \N__60534\ : std_logic;
signal \N__60531\ : std_logic;
signal \N__60528\ : std_logic;
signal \N__60523\ : std_logic;
signal \N__60522\ : std_logic;
signal \N__60521\ : std_logic;
signal \N__60520\ : std_logic;
signal \N__60519\ : std_logic;
signal \N__60518\ : std_logic;
signal \N__60517\ : std_logic;
signal \N__60516\ : std_logic;
signal \N__60513\ : std_logic;
signal \N__60510\ : std_logic;
signal \N__60507\ : std_logic;
signal \N__60502\ : std_logic;
signal \N__60501\ : std_logic;
signal \N__60500\ : std_logic;
signal \N__60499\ : std_logic;
signal \N__60498\ : std_logic;
signal \N__60497\ : std_logic;
signal \N__60496\ : std_logic;
signal \N__60495\ : std_logic;
signal \N__60490\ : std_logic;
signal \N__60487\ : std_logic;
signal \N__60480\ : std_logic;
signal \N__60479\ : std_logic;
signal \N__60478\ : std_logic;
signal \N__60475\ : std_logic;
signal \N__60470\ : std_logic;
signal \N__60469\ : std_logic;
signal \N__60468\ : std_logic;
signal \N__60467\ : std_logic;
signal \N__60464\ : std_logic;
signal \N__60463\ : std_logic;
signal \N__60462\ : std_logic;
signal \N__60461\ : std_logic;
signal \N__60458\ : std_logic;
signal \N__60453\ : std_logic;
signal \N__60446\ : std_logic;
signal \N__60439\ : std_logic;
signal \N__60436\ : std_logic;
signal \N__60433\ : std_logic;
signal \N__60426\ : std_logic;
signal \N__60423\ : std_logic;
signal \N__60416\ : std_logic;
signal \N__60413\ : std_logic;
signal \N__60410\ : std_logic;
signal \N__60407\ : std_logic;
signal \N__60398\ : std_logic;
signal \N__60397\ : std_logic;
signal \N__60396\ : std_logic;
signal \N__60395\ : std_logic;
signal \N__60392\ : std_logic;
signal \N__60389\ : std_logic;
signal \N__60386\ : std_logic;
signal \N__60381\ : std_logic;
signal \N__60376\ : std_logic;
signal \N__60371\ : std_logic;
signal \N__60366\ : std_logic;
signal \N__60359\ : std_logic;
signal \N__60358\ : std_logic;
signal \N__60357\ : std_logic;
signal \N__60354\ : std_logic;
signal \N__60353\ : std_logic;
signal \N__60352\ : std_logic;
signal \N__60349\ : std_logic;
signal \N__60344\ : std_logic;
signal \N__60341\ : std_logic;
signal \N__60336\ : std_logic;
signal \N__60331\ : std_logic;
signal \N__60326\ : std_logic;
signal \N__60321\ : std_logic;
signal \N__60318\ : std_logic;
signal \N__60315\ : std_logic;
signal \N__60314\ : std_logic;
signal \N__60313\ : std_logic;
signal \N__60310\ : std_logic;
signal \N__60309\ : std_logic;
signal \N__60304\ : std_logic;
signal \N__60301\ : std_logic;
signal \N__60294\ : std_logic;
signal \N__60285\ : std_logic;
signal \N__60282\ : std_logic;
signal \N__60273\ : std_logic;
signal \N__60270\ : std_logic;
signal \N__60269\ : std_logic;
signal \N__60266\ : std_logic;
signal \N__60263\ : std_logic;
signal \N__60262\ : std_logic;
signal \N__60251\ : std_logic;
signal \N__60250\ : std_logic;
signal \N__60249\ : std_logic;
signal \N__60248\ : std_logic;
signal \N__60247\ : std_logic;
signal \N__60240\ : std_logic;
signal \N__60237\ : std_logic;
signal \N__60234\ : std_logic;
signal \N__60233\ : std_logic;
signal \N__60230\ : std_logic;
signal \N__60225\ : std_logic;
signal \N__60212\ : std_logic;
signal \N__60209\ : std_logic;
signal \N__60204\ : std_logic;
signal \N__60195\ : std_logic;
signal \N__60186\ : std_logic;
signal \N__60181\ : std_logic;
signal \N__60176\ : std_logic;
signal \N__60173\ : std_logic;
signal \N__60170\ : std_logic;
signal \N__60167\ : std_logic;
signal \N__60164\ : std_logic;
signal \N__60157\ : std_logic;
signal \N__60154\ : std_logic;
signal \N__60151\ : std_logic;
signal \N__60148\ : std_logic;
signal \N__60143\ : std_logic;
signal \N__60132\ : std_logic;
signal \N__60123\ : std_logic;
signal \N__60100\ : std_logic;
signal \N__60099\ : std_logic;
signal \N__60098\ : std_logic;
signal \N__60097\ : std_logic;
signal \N__60096\ : std_logic;
signal \N__60095\ : std_logic;
signal \N__60094\ : std_logic;
signal \N__60093\ : std_logic;
signal \N__60092\ : std_logic;
signal \N__60091\ : std_logic;
signal \N__60090\ : std_logic;
signal \N__60087\ : std_logic;
signal \N__60084\ : std_logic;
signal \N__60083\ : std_logic;
signal \N__60082\ : std_logic;
signal \N__60081\ : std_logic;
signal \N__60080\ : std_logic;
signal \N__60077\ : std_logic;
signal \N__60076\ : std_logic;
signal \N__60073\ : std_logic;
signal \N__60072\ : std_logic;
signal \N__60069\ : std_logic;
signal \N__60066\ : std_logic;
signal \N__60065\ : std_logic;
signal \N__60064\ : std_logic;
signal \N__60063\ : std_logic;
signal \N__60060\ : std_logic;
signal \N__60059\ : std_logic;
signal \N__60058\ : std_logic;
signal \N__60053\ : std_logic;
signal \N__60052\ : std_logic;
signal \N__60049\ : std_logic;
signal \N__60048\ : std_logic;
signal \N__60047\ : std_logic;
signal \N__60046\ : std_logic;
signal \N__60045\ : std_logic;
signal \N__60044\ : std_logic;
signal \N__60043\ : std_logic;
signal \N__60042\ : std_logic;
signal \N__60041\ : std_logic;
signal \N__60040\ : std_logic;
signal \N__60037\ : std_logic;
signal \N__60036\ : std_logic;
signal \N__60031\ : std_logic;
signal \N__60026\ : std_logic;
signal \N__60021\ : std_logic;
signal \N__60018\ : std_logic;
signal \N__60015\ : std_logic;
signal \N__60014\ : std_logic;
signal \N__60009\ : std_logic;
signal \N__60008\ : std_logic;
signal \N__60007\ : std_logic;
signal \N__60006\ : std_logic;
signal \N__60003\ : std_logic;
signal \N__60002\ : std_logic;
signal \N__60001\ : std_logic;
signal \N__60000\ : std_logic;
signal \N__59999\ : std_logic;
signal \N__59996\ : std_logic;
signal \N__59995\ : std_logic;
signal \N__59994\ : std_logic;
signal \N__59993\ : std_logic;
signal \N__59992\ : std_logic;
signal \N__59991\ : std_logic;
signal \N__59988\ : std_logic;
signal \N__59987\ : std_logic;
signal \N__59986\ : std_logic;
signal \N__59985\ : std_logic;
signal \N__59984\ : std_logic;
signal \N__59983\ : std_logic;
signal \N__59982\ : std_logic;
signal \N__59979\ : std_logic;
signal \N__59978\ : std_logic;
signal \N__59977\ : std_logic;
signal \N__59976\ : std_logic;
signal \N__59975\ : std_logic;
signal \N__59974\ : std_logic;
signal \N__59973\ : std_logic;
signal \N__59970\ : std_logic;
signal \N__59969\ : std_logic;
signal \N__59966\ : std_logic;
signal \N__59965\ : std_logic;
signal \N__59964\ : std_logic;
signal \N__59963\ : std_logic;
signal \N__59962\ : std_logic;
signal \N__59961\ : std_logic;
signal \N__59960\ : std_logic;
signal \N__59955\ : std_logic;
signal \N__59954\ : std_logic;
signal \N__59951\ : std_logic;
signal \N__59944\ : std_logic;
signal \N__59937\ : std_logic;
signal \N__59936\ : std_logic;
signal \N__59933\ : std_logic;
signal \N__59930\ : std_logic;
signal \N__59925\ : std_logic;
signal \N__59922\ : std_logic;
signal \N__59917\ : std_logic;
signal \N__59912\ : std_logic;
signal \N__59905\ : std_logic;
signal \N__59904\ : std_logic;
signal \N__59901\ : std_logic;
signal \N__59900\ : std_logic;
signal \N__59897\ : std_logic;
signal \N__59894\ : std_logic;
signal \N__59891\ : std_logic;
signal \N__59888\ : std_logic;
signal \N__59887\ : std_logic;
signal \N__59884\ : std_logic;
signal \N__59881\ : std_logic;
signal \N__59874\ : std_logic;
signal \N__59871\ : std_logic;
signal \N__59868\ : std_logic;
signal \N__59867\ : std_logic;
signal \N__59862\ : std_logic;
signal \N__59857\ : std_logic;
signal \N__59854\ : std_logic;
signal \N__59851\ : std_logic;
signal \N__59846\ : std_logic;
signal \N__59839\ : std_logic;
signal \N__59836\ : std_logic;
signal \N__59831\ : std_logic;
signal \N__59828\ : std_logic;
signal \N__59823\ : std_logic;
signal \N__59822\ : std_logic;
signal \N__59819\ : std_logic;
signal \N__59816\ : std_logic;
signal \N__59813\ : std_logic;
signal \N__59812\ : std_logic;
signal \N__59809\ : std_logic;
signal \N__59802\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59785\ : std_logic;
signal \N__59780\ : std_logic;
signal \N__59777\ : std_logic;
signal \N__59772\ : std_logic;
signal \N__59769\ : std_logic;
signal \N__59764\ : std_logic;
signal \N__59759\ : std_logic;
signal \N__59756\ : std_logic;
signal \N__59751\ : std_logic;
signal \N__59748\ : std_logic;
signal \N__59743\ : std_logic;
signal \N__59740\ : std_logic;
signal \N__59737\ : std_logic;
signal \N__59734\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59722\ : std_logic;
signal \N__59717\ : std_logic;
signal \N__59704\ : std_logic;
signal \N__59703\ : std_logic;
signal \N__59702\ : std_logic;
signal \N__59697\ : std_logic;
signal \N__59692\ : std_logic;
signal \N__59687\ : std_logic;
signal \N__59684\ : std_logic;
signal \N__59673\ : std_logic;
signal \N__59672\ : std_logic;
signal \N__59661\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59649\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59629\ : std_logic;
signal \N__59624\ : std_logic;
signal \N__59619\ : std_logic;
signal \N__59612\ : std_logic;
signal \N__59609\ : std_logic;
signal \N__59606\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59584\ : std_logic;
signal \N__59581\ : std_logic;
signal \N__59578\ : std_logic;
signal \N__59575\ : std_logic;
signal \N__59572\ : std_logic;
signal \N__59569\ : std_logic;
signal \N__59566\ : std_logic;
signal \N__59563\ : std_logic;
signal \N__59560\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59551\ : std_logic;
signal \N__59548\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59542\ : std_logic;
signal \N__59539\ : std_logic;
signal \N__59536\ : std_logic;
signal \N__59533\ : std_logic;
signal \N__59530\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59524\ : std_logic;
signal \N__59521\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59516\ : std_logic;
signal \N__59515\ : std_logic;
signal \N__59514\ : std_logic;
signal \N__59513\ : std_logic;
signal \N__59510\ : std_logic;
signal \N__59509\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59507\ : std_logic;
signal \N__59506\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59504\ : std_logic;
signal \N__59503\ : std_logic;
signal \N__59502\ : std_logic;
signal \N__59501\ : std_logic;
signal \N__59498\ : std_logic;
signal \N__59497\ : std_logic;
signal \N__59496\ : std_logic;
signal \N__59493\ : std_logic;
signal \N__59492\ : std_logic;
signal \N__59491\ : std_logic;
signal \N__59490\ : std_logic;
signal \N__59489\ : std_logic;
signal \N__59488\ : std_logic;
signal \N__59485\ : std_logic;
signal \N__59484\ : std_logic;
signal \N__59483\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59479\ : std_logic;
signal \N__59476\ : std_logic;
signal \N__59475\ : std_logic;
signal \N__59472\ : std_logic;
signal \N__59469\ : std_logic;
signal \N__59468\ : std_logic;
signal \N__59467\ : std_logic;
signal \N__59466\ : std_logic;
signal \N__59461\ : std_logic;
signal \N__59458\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59450\ : std_logic;
signal \N__59447\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59444\ : std_logic;
signal \N__59443\ : std_logic;
signal \N__59442\ : std_logic;
signal \N__59441\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59439\ : std_logic;
signal \N__59438\ : std_logic;
signal \N__59437\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59435\ : std_logic;
signal \N__59434\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59432\ : std_logic;
signal \N__59431\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59429\ : std_logic;
signal \N__59428\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59425\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59423\ : std_logic;
signal \N__59422\ : std_logic;
signal \N__59421\ : std_logic;
signal \N__59420\ : std_logic;
signal \N__59417\ : std_logic;
signal \N__59414\ : std_logic;
signal \N__59411\ : std_logic;
signal \N__59410\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59408\ : std_logic;
signal \N__59407\ : std_logic;
signal \N__59406\ : std_logic;
signal \N__59405\ : std_logic;
signal \N__59402\ : std_logic;
signal \N__59401\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59399\ : std_logic;
signal \N__59398\ : std_logic;
signal \N__59397\ : std_logic;
signal \N__59394\ : std_logic;
signal \N__59391\ : std_logic;
signal \N__59388\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59378\ : std_logic;
signal \N__59373\ : std_logic;
signal \N__59372\ : std_logic;
signal \N__59371\ : std_logic;
signal \N__59368\ : std_logic;
signal \N__59367\ : std_logic;
signal \N__59366\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59364\ : std_logic;
signal \N__59363\ : std_logic;
signal \N__59362\ : std_logic;
signal \N__59359\ : std_logic;
signal \N__59356\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59354\ : std_logic;
signal \N__59353\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59351\ : std_logic;
signal \N__59350\ : std_logic;
signal \N__59347\ : std_logic;
signal \N__59342\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59335\ : std_logic;
signal \N__59332\ : std_logic;
signal \N__59331\ : std_logic;
signal \N__59330\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59327\ : std_logic;
signal \N__59326\ : std_logic;
signal \N__59325\ : std_logic;
signal \N__59324\ : std_logic;
signal \N__59323\ : std_logic;
signal \N__59322\ : std_logic;
signal \N__59321\ : std_logic;
signal \N__59320\ : std_logic;
signal \N__59317\ : std_logic;
signal \N__59308\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59306\ : std_logic;
signal \N__59305\ : std_logic;
signal \N__59298\ : std_logic;
signal \N__59293\ : std_logic;
signal \N__59288\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59278\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59268\ : std_logic;
signal \N__59267\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59265\ : std_logic;
signal \N__59264\ : std_logic;
signal \N__59263\ : std_logic;
signal \N__59262\ : std_logic;
signal \N__59261\ : std_logic;
signal \N__59258\ : std_logic;
signal \N__59251\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59246\ : std_logic;
signal \N__59241\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59231\ : std_logic;
signal \N__59228\ : std_logic;
signal \N__59227\ : std_logic;
signal \N__59226\ : std_logic;
signal \N__59225\ : std_logic;
signal \N__59218\ : std_logic;
signal \N__59215\ : std_logic;
signal \N__59210\ : std_logic;
signal \N__59209\ : std_logic;
signal \N__59206\ : std_logic;
signal \N__59201\ : std_logic;
signal \N__59198\ : std_logic;
signal \N__59193\ : std_logic;
signal \N__59192\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59189\ : std_logic;
signal \N__59186\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59182\ : std_logic;
signal \N__59181\ : std_logic;
signal \N__59178\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59160\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59127\ : std_logic;
signal \N__59124\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59116\ : std_logic;
signal \N__59115\ : std_logic;
signal \N__59114\ : std_logic;
signal \N__59113\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59106\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59094\ : std_logic;
signal \N__59091\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59079\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__59069\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59063\ : std_logic;
signal \N__59060\ : std_logic;
signal \N__59057\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59045\ : std_logic;
signal \N__59042\ : std_logic;
signal \N__59035\ : std_logic;
signal \N__59026\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59020\ : std_logic;
signal \N__59017\ : std_logic;
signal \N__59016\ : std_logic;
signal \N__59015\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59010\ : std_logic;
signal \N__59009\ : std_logic;
signal \N__59006\ : std_logic;
signal \N__58999\ : std_logic;
signal \N__58996\ : std_logic;
signal \N__58993\ : std_logic;
signal \N__58988\ : std_logic;
signal \N__58981\ : std_logic;
signal \N__58978\ : std_logic;
signal \N__58973\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58963\ : std_logic;
signal \N__58960\ : std_logic;
signal \N__58957\ : std_logic;
signal \N__58954\ : std_logic;
signal \N__58951\ : std_logic;
signal \N__58950\ : std_logic;
signal \N__58949\ : std_logic;
signal \N__58948\ : std_logic;
signal \N__58945\ : std_logic;
signal \N__58942\ : std_logic;
signal \N__58939\ : std_logic;
signal \N__58934\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58916\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58908\ : std_logic;
signal \N__58905\ : std_logic;
signal \N__58902\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58889\ : std_logic;
signal \N__58870\ : std_logic;
signal \N__58861\ : std_logic;
signal \N__58858\ : std_logic;
signal \N__58857\ : std_logic;
signal \N__58856\ : std_logic;
signal \N__58855\ : std_logic;
signal \N__58852\ : std_logic;
signal \N__58845\ : std_logic;
signal \N__58844\ : std_logic;
signal \N__58843\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58841\ : std_logic;
signal \N__58840\ : std_logic;
signal \N__58837\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58831\ : std_logic;
signal \N__58828\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58814\ : std_logic;
signal \N__58807\ : std_logic;
signal \N__58798\ : std_logic;
signal \N__58791\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58777\ : std_logic;
signal \N__58774\ : std_logic;
signal \N__58771\ : std_logic;
signal \N__58766\ : std_logic;
signal \N__58753\ : std_logic;
signal \N__58746\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58740\ : std_logic;
signal \N__58733\ : std_logic;
signal \N__58730\ : std_logic;
signal \N__58727\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58721\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58700\ : std_logic;
signal \N__58689\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58654\ : std_logic;
signal \N__58653\ : std_logic;
signal \N__58652\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58650\ : std_logic;
signal \N__58649\ : std_logic;
signal \N__58648\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58642\ : std_logic;
signal \N__58641\ : std_logic;
signal \N__58638\ : std_logic;
signal \N__58635\ : std_logic;
signal \N__58630\ : std_logic;
signal \N__58627\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58625\ : std_logic;
signal \N__58624\ : std_logic;
signal \N__58621\ : std_logic;
signal \N__58616\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58614\ : std_logic;
signal \N__58611\ : std_logic;
signal \N__58610\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58608\ : std_logic;
signal \N__58607\ : std_logic;
signal \N__58602\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58594\ : std_logic;
signal \N__58591\ : std_logic;
signal \N__58586\ : std_logic;
signal \N__58585\ : std_logic;
signal \N__58584\ : std_logic;
signal \N__58581\ : std_logic;
signal \N__58578\ : std_logic;
signal \N__58575\ : std_logic;
signal \N__58572\ : std_logic;
signal \N__58567\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58557\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58547\ : std_logic;
signal \N__58528\ : std_logic;
signal \N__58527\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58523\ : std_logic;
signal \N__58522\ : std_logic;
signal \N__58521\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58515\ : std_logic;
signal \N__58512\ : std_logic;
signal \N__58511\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58505\ : std_logic;
signal \N__58502\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58496\ : std_logic;
signal \N__58493\ : std_logic;
signal \N__58492\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58488\ : std_logic;
signal \N__58487\ : std_logic;
signal \N__58484\ : std_logic;
signal \N__58483\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58475\ : std_logic;
signal \N__58470\ : std_logic;
signal \N__58469\ : std_logic;
signal \N__58466\ : std_logic;
signal \N__58463\ : std_logic;
signal \N__58460\ : std_logic;
signal \N__58457\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58447\ : std_logic;
signal \N__58442\ : std_logic;
signal \N__58429\ : std_logic;
signal \N__58426\ : std_logic;
signal \N__58423\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58414\ : std_logic;
signal \N__58411\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58407\ : std_logic;
signal \N__58404\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58393\ : std_logic;
signal \N__58390\ : std_logic;
signal \N__58387\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58375\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58369\ : std_logic;
signal \N__58366\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58348\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58342\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58333\ : std_logic;
signal \N__58330\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58315\ : std_logic;
signal \N__58312\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58306\ : std_logic;
signal \N__58303\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58297\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58285\ : std_logic;
signal \N__58282\ : std_logic;
signal \N__58279\ : std_logic;
signal \N__58276\ : std_logic;
signal \N__58273\ : std_logic;
signal \N__58270\ : std_logic;
signal \N__58267\ : std_logic;
signal \N__58264\ : std_logic;
signal \N__58261\ : std_logic;
signal \N__58258\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58249\ : std_logic;
signal \N__58246\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58240\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58234\ : std_logic;
signal \N__58231\ : std_logic;
signal \N__58228\ : std_logic;
signal \N__58225\ : std_logic;
signal \N__58222\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58213\ : std_logic;
signal \N__58210\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58208\ : std_logic;
signal \N__58207\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58205\ : std_logic;
signal \N__58204\ : std_logic;
signal \N__58201\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58192\ : std_logic;
signal \N__58189\ : std_logic;
signal \N__58188\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58185\ : std_logic;
signal \N__58182\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58178\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58170\ : std_logic;
signal \N__58161\ : std_logic;
signal \N__58154\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58152\ : std_logic;
signal \N__58151\ : std_logic;
signal \N__58148\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58144\ : std_logic;
signal \N__58141\ : std_logic;
signal \N__58138\ : std_logic;
signal \N__58133\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58126\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58118\ : std_logic;
signal \N__58117\ : std_logic;
signal \N__58114\ : std_logic;
signal \N__58107\ : std_logic;
signal \N__58104\ : std_logic;
signal \N__58097\ : std_logic;
signal \N__58092\ : std_logic;
signal \N__58089\ : std_logic;
signal \N__58086\ : std_logic;
signal \N__58083\ : std_logic;
signal \N__58080\ : std_logic;
signal \N__58077\ : std_logic;
signal \N__58074\ : std_logic;
signal \N__58071\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58063\ : std_logic;
signal \N__58060\ : std_logic;
signal \N__58055\ : std_logic;
signal \N__58052\ : std_logic;
signal \N__58047\ : std_logic;
signal \N__58042\ : std_logic;
signal \N__58041\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58039\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58037\ : std_logic;
signal \N__58036\ : std_logic;
signal \N__58035\ : std_logic;
signal \N__58034\ : std_logic;
signal \N__58033\ : std_logic;
signal \N__58032\ : std_logic;
signal \N__58031\ : std_logic;
signal \N__58030\ : std_logic;
signal \N__58023\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58019\ : std_logic;
signal \N__58018\ : std_logic;
signal \N__58011\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57999\ : std_logic;
signal \N__57996\ : std_logic;
signal \N__57993\ : std_logic;
signal \N__57990\ : std_logic;
signal \N__57985\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57961\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57954\ : std_logic;
signal \N__57953\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57947\ : std_logic;
signal \N__57942\ : std_logic;
signal \N__57937\ : std_logic;
signal \N__57934\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57928\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57919\ : std_logic;
signal \N__57916\ : std_logic;
signal \N__57913\ : std_logic;
signal \N__57910\ : std_logic;
signal \N__57907\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57892\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57883\ : std_logic;
signal \N__57880\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57873\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57870\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57864\ : std_logic;
signal \N__57863\ : std_logic;
signal \N__57862\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57857\ : std_logic;
signal \N__57856\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57854\ : std_logic;
signal \N__57853\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57851\ : std_logic;
signal \N__57850\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57848\ : std_logic;
signal \N__57845\ : std_logic;
signal \N__57844\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57838\ : std_logic;
signal \N__57835\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57821\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57811\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57805\ : std_logic;
signal \N__57802\ : std_logic;
signal \N__57799\ : std_logic;
signal \N__57794\ : std_logic;
signal \N__57789\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57783\ : std_logic;
signal \N__57780\ : std_logic;
signal \N__57779\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57775\ : std_logic;
signal \N__57772\ : std_logic;
signal \N__57765\ : std_logic;
signal \N__57764\ : std_logic;
signal \N__57763\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57757\ : std_logic;
signal \N__57754\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57748\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57746\ : std_logic;
signal \N__57745\ : std_logic;
signal \N__57742\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57739\ : std_logic;
signal \N__57736\ : std_logic;
signal \N__57731\ : std_logic;
signal \N__57730\ : std_logic;
signal \N__57729\ : std_logic;
signal \N__57728\ : std_logic;
signal \N__57723\ : std_logic;
signal \N__57716\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57712\ : std_logic;
signal \N__57711\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57709\ : std_logic;
signal \N__57708\ : std_logic;
signal \N__57707\ : std_logic;
signal \N__57706\ : std_logic;
signal \N__57705\ : std_logic;
signal \N__57704\ : std_logic;
signal \N__57703\ : std_logic;
signal \N__57702\ : std_logic;
signal \N__57701\ : std_logic;
signal \N__57700\ : std_logic;
signal \N__57697\ : std_logic;
signal \N__57694\ : std_logic;
signal \N__57693\ : std_logic;
signal \N__57692\ : std_logic;
signal \N__57687\ : std_logic;
signal \N__57684\ : std_logic;
signal \N__57681\ : std_logic;
signal \N__57678\ : std_logic;
signal \N__57673\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57665\ : std_logic;
signal \N__57662\ : std_logic;
signal \N__57661\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57647\ : std_logic;
signal \N__57644\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57625\ : std_logic;
signal \N__57622\ : std_logic;
signal \N__57621\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57618\ : std_logic;
signal \N__57617\ : std_logic;
signal \N__57614\ : std_logic;
signal \N__57611\ : std_logic;
signal \N__57610\ : std_logic;
signal \N__57607\ : std_logic;
signal \N__57604\ : std_logic;
signal \N__57603\ : std_logic;
signal \N__57600\ : std_logic;
signal \N__57591\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57587\ : std_logic;
signal \N__57584\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57566\ : std_logic;
signal \N__57563\ : std_logic;
signal \N__57560\ : std_logic;
signal \N__57557\ : std_logic;
signal \N__57554\ : std_logic;
signal \N__57551\ : std_logic;
signal \N__57546\ : std_logic;
signal \N__57543\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57527\ : std_logic;
signal \N__57522\ : std_logic;
signal \N__57521\ : std_logic;
signal \N__57520\ : std_logic;
signal \N__57517\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57509\ : std_logic;
signal \N__57506\ : std_logic;
signal \N__57501\ : std_logic;
signal \N__57498\ : std_logic;
signal \N__57489\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57475\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57468\ : std_logic;
signal \N__57465\ : std_logic;
signal \N__57462\ : std_logic;
signal \N__57455\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57445\ : std_logic;
signal \N__57438\ : std_logic;
signal \N__57435\ : std_logic;
signal \N__57432\ : std_logic;
signal \N__57429\ : std_logic;
signal \N__57408\ : std_logic;
signal \N__57405\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57397\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57380\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57364\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57358\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57354\ : std_logic;
signal \N__57353\ : std_logic;
signal \N__57350\ : std_logic;
signal \N__57347\ : std_logic;
signal \N__57344\ : std_logic;
signal \N__57337\ : std_logic;
signal \N__57334\ : std_logic;
signal \N__57331\ : std_logic;
signal \N__57328\ : std_logic;
signal \N__57325\ : std_logic;
signal \N__57322\ : std_logic;
signal \N__57319\ : std_logic;
signal \N__57316\ : std_logic;
signal \N__57313\ : std_logic;
signal \N__57310\ : std_logic;
signal \N__57307\ : std_logic;
signal \N__57304\ : std_logic;
signal \N__57301\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57299\ : std_logic;
signal \N__57296\ : std_logic;
signal \N__57293\ : std_logic;
signal \N__57290\ : std_logic;
signal \N__57283\ : std_logic;
signal \N__57280\ : std_logic;
signal \N__57277\ : std_logic;
signal \N__57274\ : std_logic;
signal \N__57271\ : std_logic;
signal \N__57268\ : std_logic;
signal \N__57265\ : std_logic;
signal \N__57262\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57255\ : std_logic;
signal \N__57252\ : std_logic;
signal \N__57249\ : std_logic;
signal \N__57244\ : std_logic;
signal \N__57243\ : std_logic;
signal \N__57240\ : std_logic;
signal \N__57237\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57231\ : std_logic;
signal \N__57228\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57222\ : std_logic;
signal \N__57217\ : std_logic;
signal \N__57216\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57210\ : std_logic;
signal \N__57205\ : std_logic;
signal \N__57202\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57195\ : std_logic;
signal \N__57192\ : std_logic;
signal \N__57189\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57183\ : std_logic;
signal \N__57178\ : std_logic;
signal \N__57177\ : std_logic;
signal \N__57176\ : std_logic;
signal \N__57175\ : std_logic;
signal \N__57174\ : std_logic;
signal \N__57173\ : std_logic;
signal \N__57172\ : std_logic;
signal \N__57171\ : std_logic;
signal \N__57170\ : std_logic;
signal \N__57167\ : std_logic;
signal \N__57164\ : std_logic;
signal \N__57161\ : std_logic;
signal \N__57148\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57138\ : std_logic;
signal \N__57137\ : std_logic;
signal \N__57136\ : std_logic;
signal \N__57135\ : std_logic;
signal \N__57132\ : std_logic;
signal \N__57131\ : std_logic;
signal \N__57130\ : std_logic;
signal \N__57129\ : std_logic;
signal \N__57126\ : std_logic;
signal \N__57123\ : std_logic;
signal \N__57122\ : std_logic;
signal \N__57121\ : std_logic;
signal \N__57120\ : std_logic;
signal \N__57119\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57117\ : std_logic;
signal \N__57116\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57113\ : std_logic;
signal \N__57112\ : std_logic;
signal \N__57111\ : std_logic;
signal \N__57110\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57100\ : std_logic;
signal \N__57097\ : std_logic;
signal \N__57096\ : std_logic;
signal \N__57093\ : std_logic;
signal \N__57092\ : std_logic;
signal \N__57087\ : std_logic;
signal \N__57084\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57078\ : std_logic;
signal \N__57077\ : std_logic;
signal \N__57074\ : std_logic;
signal \N__57071\ : std_logic;
signal \N__57070\ : std_logic;
signal \N__57063\ : std_logic;
signal \N__57058\ : std_logic;
signal \N__57053\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57049\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57037\ : std_logic;
signal \N__57034\ : std_logic;
signal \N__57031\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57022\ : std_logic;
signal \N__57019\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57011\ : std_logic;
signal \N__57008\ : std_logic;
signal \N__57003\ : std_logic;
signal \N__57000\ : std_logic;
signal \N__56997\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56989\ : std_logic;
signal \N__56984\ : std_logic;
signal \N__56979\ : std_logic;
signal \N__56972\ : std_logic;
signal \N__56969\ : std_logic;
signal \N__56962\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56950\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56933\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56923\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56908\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56896\ : std_logic;
signal \N__56893\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56887\ : std_logic;
signal \N__56884\ : std_logic;
signal \N__56881\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56872\ : std_logic;
signal \N__56871\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56862\ : std_logic;
signal \N__56859\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56851\ : std_logic;
signal \N__56850\ : std_logic;
signal \N__56849\ : std_logic;
signal \N__56846\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56840\ : std_logic;
signal \N__56839\ : std_logic;
signal \N__56838\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56831\ : std_logic;
signal \N__56828\ : std_logic;
signal \N__56825\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56819\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56813\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56793\ : std_logic;
signal \N__56790\ : std_logic;
signal \N__56785\ : std_logic;
signal \N__56776\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56770\ : std_logic;
signal \N__56767\ : std_logic;
signal \N__56764\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56740\ : std_logic;
signal \N__56739\ : std_logic;
signal \N__56736\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56730\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56722\ : std_logic;
signal \N__56721\ : std_logic;
signal \N__56718\ : std_logic;
signal \N__56715\ : std_logic;
signal \N__56710\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56706\ : std_logic;
signal \N__56703\ : std_logic;
signal \N__56700\ : std_logic;
signal \N__56697\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56689\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56685\ : std_logic;
signal \N__56682\ : std_logic;
signal \N__56677\ : std_logic;
signal \N__56676\ : std_logic;
signal \N__56673\ : std_logic;
signal \N__56670\ : std_logic;
signal \N__56667\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56658\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56647\ : std_logic;
signal \N__56644\ : std_logic;
signal \N__56643\ : std_logic;
signal \N__56640\ : std_logic;
signal \N__56637\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56628\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56622\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56613\ : std_logic;
signal \N__56610\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56602\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56592\ : std_logic;
signal \N__56587\ : std_logic;
signal \N__56584\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56577\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56570\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56566\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56548\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56540\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56532\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56503\ : std_logic;
signal \N__56502\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56496\ : std_logic;
signal \N__56495\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56475\ : std_logic;
signal \N__56474\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56470\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56463\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56460\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56458\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56439\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56429\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56423\ : std_logic;
signal \N__56420\ : std_logic;
signal \N__56417\ : std_logic;
signal \N__56414\ : std_logic;
signal \N__56405\ : std_logic;
signal \N__56396\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56386\ : std_logic;
signal \N__56383\ : std_logic;
signal \N__56380\ : std_logic;
signal \N__56377\ : std_logic;
signal \N__56376\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56365\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56356\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56350\ : std_logic;
signal \N__56347\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56332\ : std_logic;
signal \N__56329\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56310\ : std_logic;
signal \N__56307\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56274\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56222\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56212\ : std_logic;
signal \N__56209\ : std_logic;
signal \N__56206\ : std_logic;
signal \N__56205\ : std_logic;
signal \N__56202\ : std_logic;
signal \N__56199\ : std_logic;
signal \N__56196\ : std_logic;
signal \N__56193\ : std_logic;
signal \N__56190\ : std_logic;
signal \N__56185\ : std_logic;
signal \N__56184\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56178\ : std_logic;
signal \N__56173\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56167\ : std_logic;
signal \N__56164\ : std_logic;
signal \N__56161\ : std_logic;
signal \N__56158\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56142\ : std_logic;
signal \N__56137\ : std_logic;
signal \N__56134\ : std_logic;
signal \N__56133\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56123\ : std_logic;
signal \N__56120\ : std_logic;
signal \N__56117\ : std_logic;
signal \N__56110\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56078\ : std_logic;
signal \N__56075\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56066\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56045\ : std_logic;
signal \N__56042\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56023\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56019\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56004\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55987\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55963\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55954\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55948\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55942\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55936\ : std_logic;
signal \N__55935\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55925\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55914\ : std_logic;
signal \N__55909\ : std_logic;
signal \N__55906\ : std_logic;
signal \N__55903\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55896\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55881\ : std_logic;
signal \N__55878\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55870\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55852\ : std_logic;
signal \N__55849\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55845\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55841\ : std_logic;
signal \N__55838\ : std_logic;
signal \N__55837\ : std_logic;
signal \N__55834\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55828\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55822\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55802\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55784\ : std_logic;
signal \N__55781\ : std_logic;
signal \N__55774\ : std_logic;
signal \N__55771\ : std_logic;
signal \N__55770\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55764\ : std_logic;
signal \N__55761\ : std_logic;
signal \N__55758\ : std_logic;
signal \N__55755\ : std_logic;
signal \N__55752\ : std_logic;
signal \N__55751\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55721\ : std_logic;
signal \N__55714\ : std_logic;
signal \N__55711\ : std_logic;
signal \N__55710\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55708\ : std_logic;
signal \N__55707\ : std_logic;
signal \N__55704\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55700\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55691\ : std_logic;
signal \N__55686\ : std_logic;
signal \N__55683\ : std_logic;
signal \N__55678\ : std_logic;
signal \N__55675\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55658\ : std_logic;
signal \N__55651\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55649\ : std_logic;
signal \N__55646\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55640\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55636\ : std_logic;
signal \N__55635\ : std_logic;
signal \N__55634\ : std_logic;
signal \N__55631\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55616\ : std_logic;
signal \N__55613\ : std_logic;
signal \N__55610\ : std_logic;
signal \N__55607\ : std_logic;
signal \N__55604\ : std_logic;
signal \N__55599\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55576\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55570\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55542\ : std_logic;
signal \N__55539\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55529\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55520\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55498\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55487\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55474\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55461\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55401\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55394\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55385\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55380\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55372\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55369\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55338\ : std_logic;
signal \N__55335\ : std_logic;
signal \N__55332\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55323\ : std_logic;
signal \N__55320\ : std_logic;
signal \N__55313\ : std_logic;
signal \N__55310\ : std_logic;
signal \N__55307\ : std_logic;
signal \N__55304\ : std_logic;
signal \N__55297\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55277\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55267\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55261\ : std_logic;
signal \N__55258\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55249\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55203\ : std_logic;
signal \N__55200\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55194\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55170\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55139\ : std_logic;
signal \N__55136\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55099\ : std_logic;
signal \N__55096\ : std_logic;
signal \N__55093\ : std_logic;
signal \N__55090\ : std_logic;
signal \N__55087\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55081\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55072\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55051\ : std_logic;
signal \N__55048\ : std_logic;
signal \N__55045\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55039\ : std_logic;
signal \N__55038\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55025\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55016\ : std_logic;
signal \N__55013\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55003\ : std_logic;
signal \N__55000\ : std_logic;
signal \N__54991\ : std_logic;
signal \N__54988\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54982\ : std_logic;
signal \N__54979\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54970\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54964\ : std_logic;
signal \N__54961\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54949\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54943\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54939\ : std_logic;
signal \N__54938\ : std_logic;
signal \N__54935\ : std_logic;
signal \N__54932\ : std_logic;
signal \N__54931\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54926\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54920\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54897\ : std_logic;
signal \N__54896\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54850\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54826\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54820\ : std_logic;
signal \N__54817\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54809\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54801\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54797\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54793\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54782\ : std_logic;
signal \N__54779\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54769\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54735\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54712\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54682\ : std_logic;
signal \N__54679\ : std_logic;
signal \N__54676\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54666\ : std_logic;
signal \N__54663\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54651\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54647\ : std_logic;
signal \N__54644\ : std_logic;
signal \N__54641\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54622\ : std_logic;
signal \N__54619\ : std_logic;
signal \N__54616\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54608\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54602\ : std_logic;
signal \N__54601\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54587\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54578\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54572\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54562\ : std_logic;
signal \N__54559\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54542\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54539\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54537\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54529\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54527\ : std_logic;
signal \N__54526\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54487\ : std_logic;
signal \N__54484\ : std_logic;
signal \N__54475\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54465\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54445\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54430\ : std_logic;
signal \N__54427\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54415\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54409\ : std_logic;
signal \N__54408\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54391\ : std_logic;
signal \N__54388\ : std_logic;
signal \N__54385\ : std_logic;
signal \N__54382\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54372\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54353\ : std_logic;
signal \N__54350\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54330\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54313\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54311\ : std_logic;
signal \N__54310\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54307\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54282\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54264\ : std_logic;
signal \N__54259\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54234\ : std_logic;
signal \N__54231\ : std_logic;
signal \N__54220\ : std_logic;
signal \N__54205\ : std_logic;
signal \N__54202\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54195\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54189\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54182\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54171\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54162\ : std_logic;
signal \N__54161\ : std_logic;
signal \N__54160\ : std_logic;
signal \N__54159\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54153\ : std_logic;
signal \N__54150\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54137\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54125\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54116\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54110\ : std_logic;
signal \N__54101\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54072\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54065\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54049\ : std_logic;
signal \N__54044\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54017\ : std_logic;
signal \N__54016\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53935\ : std_logic;
signal \N__53932\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53923\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53914\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53896\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53893\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53857\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53855\ : std_logic;
signal \N__53852\ : std_logic;
signal \N__53847\ : std_logic;
signal \N__53844\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53824\ : std_logic;
signal \N__53821\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53800\ : std_logic;
signal \N__53797\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53781\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53739\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53736\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53733\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53707\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53703\ : std_logic;
signal \N__53700\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53692\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53678\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53671\ : std_logic;
signal \N__53670\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53665\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53653\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53638\ : std_logic;
signal \N__53635\ : std_logic;
signal \N__53634\ : std_logic;
signal \N__53631\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53624\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53617\ : std_logic;
signal \N__53614\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53606\ : std_logic;
signal \N__53603\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53598\ : std_logic;
signal \N__53595\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53588\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53580\ : std_logic;
signal \N__53577\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53569\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53558\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53504\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53473\ : std_logic;
signal \N__53464\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53443\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53432\ : std_logic;
signal \N__53429\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53416\ : std_logic;
signal \N__53413\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53391\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53361\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53353\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53338\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53314\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53307\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53301\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53287\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53233\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53197\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53191\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53182\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53164\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53148\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53107\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53101\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53083\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53049\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53035\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53026\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52926\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52913\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52909\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52850\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52842\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52829\ : std_logic;
signal \N__52826\ : std_logic;
signal \N__52823\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52805\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52783\ : std_logic;
signal \N__52780\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52733\ : std_logic;
signal \N__52730\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52717\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52681\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52658\ : std_logic;
signal \N__52655\ : std_logic;
signal \N__52652\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52642\ : std_logic;
signal \N__52639\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52622\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52575\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52502\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52273\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52193\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52142\ : std_logic;
signal \N__52139\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52115\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52101\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51965\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51941\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51831\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51615\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51560\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51546\ : std_logic;
signal \N__51543\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51459\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51354\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51141\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51052\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51036\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51028\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51007\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50998\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50862\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50738\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50627\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\ : std_logic;
signal \RTD_SCLK\ : std_logic;
signal \RTD.n8\ : std_logic;
signal \RTD_SDI\ : std_logic;
signal \RTD.n21253\ : std_logic;
signal \VAC_MISO\ : std_logic;
signal cmd_rdadctmp_0_adj_1548 : std_logic;
signal \VAC_SCLK\ : std_logic;
signal \n14_cascade_\ : std_logic;
signal n21889 : std_logic;
signal \VAC_CS\ : std_logic;
signal \DDS_SCK1\ : std_logic;
signal \RTD.n12262\ : std_logic;
signal \RTD_SDO\ : std_logic;
signal \CLK_DDS.n18366\ : std_logic;
signal bit_cnt_0_adj_1512 : std_logic;
signal bit_cnt_3 : std_logic;
signal n22326 : std_logic;
signal \CLK_DDS.n9\ : std_logic;
signal buf_adcdata_vac_4 : std_logic;
signal cmd_rdadctmp_1_adj_1547 : std_logic;
signal cmd_rdadctmp_14_adj_1534 : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \ADC_VAC.n20683\ : std_logic;
signal \ADC_VAC.n20684\ : std_logic;
signal \ADC_VAC.n20685\ : std_logic;
signal \ADC_VAC.n20686\ : std_logic;
signal \ADC_VAC.n20687\ : std_logic;
signal \ADC_VAC.n20688\ : std_logic;
signal \ADC_VAC.n20689\ : std_logic;
signal \ADC_VAC.n13784\ : std_logic;
signal \ADC_VAC.n13784_cascade_\ : std_logic;
signal \ADC_VAC.n15660\ : std_logic;
signal \RTD.n22632_cascade_\ : std_logic;
signal \DDS_CS1\ : std_logic;
signal \CLK_DDS.n9_adj_1489\ : std_logic;
signal read_buf_15 : std_logic;
signal read_buf_10 : std_logic;
signal bit_cnt_2 : std_logic;
signal bit_cnt_1 : std_logic;
signal dds_state_0_adj_1510 : std_logic;
signal n8_adj_1686 : std_logic;
signal read_buf_11 : std_logic;
signal read_buf_12 : std_logic;
signal read_buf_14 : std_logic;
signal read_buf_3 : std_logic;
signal read_buf_13 : std_logic;
signal \n19_adj_1690_cascade_\ : std_logic;
signal buf_adcdata_vac_6 : std_logic;
signal \n19_adj_1693_cascade_\ : std_logic;
signal buf_data_iac_5 : std_logic;
signal buf_adcdata_iac_6 : std_logic;
signal buf_adcdata_iac_7 : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal n19_adj_1700 : std_logic;
signal buf_data_iac_4 : std_logic;
signal \n22_adj_1701_cascade_\ : std_logic;
signal buf_adcdata_vac_7 : std_logic;
signal buf_adcdata_iac_4 : std_logic;
signal n22_adj_1697 : std_logic;
signal cmd_rdadctmp_15_adj_1533 : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal buf_adcdata_iac_5 : std_logic;
signal \ADC_VAC.n13747_cascade_\ : std_logic;
signal \ADC_VAC.n13842\ : std_logic;
signal \ADC_VAC.bit_cnt_2\ : std_logic;
signal \ADC_VAC.bit_cnt_1\ : std_logic;
signal \ADC_VAC.bit_cnt_3\ : std_logic;
signal \ADC_VAC.bit_cnt_4\ : std_logic;
signal \ADC_VAC.bit_cnt_6\ : std_logic;
signal \ADC_VAC.bit_cnt_0\ : std_logic;
signal \ADC_VAC.n22109_cascade_\ : std_logic;
signal \ADC_VAC.bit_cnt_7\ : std_logic;
signal \ADC_VAC.n22126_cascade_\ : std_logic;
signal \ADC_VAC.bit_cnt_5\ : std_logic;
signal \ADC_VAC.n22389_cascade_\ : std_logic;
signal \ADC_VAC.n22030\ : std_logic;
signal \ADC_VAC.n17\ : std_logic;
signal \VAC_DRDY\ : std_logic;
signal \ADC_VAC.n12\ : std_logic;
signal \RTD_CS\ : std_logic;
signal \RTD.n22382\ : std_logic;
signal \RTD.n20051_cascade_\ : std_logic;
signal \RTD.n22079\ : std_logic;
signal \RTD.n22599_cascade_\ : std_logic;
signal \RTD.n23689\ : std_logic;
signal \RTD.n56_cascade_\ : std_logic;
signal \RTD.n5\ : std_logic;
signal \RTD.n71\ : std_logic;
signal \RTD.n71_cascade_\ : std_logic;
signal \RTD.n22623\ : std_logic;
signal \RTD.n20051\ : std_logic;
signal read_buf_0 : std_logic;
signal \RTD.read_buf_4\ : std_logic;
signal \n21989_cascade_\ : std_logic;
signal read_buf_1 : std_logic;
signal read_buf_2 : std_logic;
signal \RTD.n68_cascade_\ : std_logic;
signal \RTD.cfg_buf_4\ : std_logic;
signal \RTD.cfg_buf_2\ : std_logic;
signal \RTD.cfg_buf_0\ : std_logic;
signal \RTD.n10\ : std_logic;
signal \RTD.n9_cascade_\ : std_logic;
signal \RTD.cfg_buf_3\ : std_logic;
signal \RTD.adress_7\ : std_logic;
signal \RTD.n19_cascade_\ : std_logic;
signal \RTD.n15396\ : std_logic;
signal \RTD.n1\ : std_logic;
signal \RTD.n1_cascade_\ : std_logic;
signal \RTD.cfg_tmp_0\ : std_logic;
signal \RTD.cfg_tmp_1\ : std_logic;
signal \RTD.cfg_tmp_2\ : std_logic;
signal \RTD.cfg_tmp_3\ : std_logic;
signal \RTD.cfg_tmp_4\ : std_logic;
signal \RTD.cfg_tmp_5\ : std_logic;
signal \RTD.cfg_tmp_6\ : std_logic;
signal \RTD.cfg_tmp_7\ : std_logic;
signal buf_data_iac_6 : std_logic;
signal n22_adj_1694 : std_logic;
signal \buf_readRTD_1\ : std_logic;
signal cmd_rdadctmp_2_adj_1546 : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal n19_adj_1696 : std_logic;
signal buf_data_iac_7 : std_logic;
signal n22_adj_1691 : std_logic;
signal cmd_rdadctmp_16_adj_1532 : std_logic;
signal cmd_rdadctmp_23_adj_1525 : std_logic;
signal cmd_rdadctmp_24_adj_1524 : std_logic;
signal cmd_rdadctmp_28_adj_1520 : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal cmd_rdadctmp_13_adj_1535 : std_logic;
signal buf_adcdata_vac_5 : std_logic;
signal cmd_rdadctmp_17_adj_1531 : std_logic;
signal cmd_rdadctmp_18_adj_1530 : std_logic;
signal \n23543_cascade_\ : std_logic;
signal cmd_rdadctmp_31_adj_1517 : std_logic;
signal cmd_rdadctmp_29_adj_1519 : std_logic;
signal cmd_rdadctmp_30_adj_1518 : std_logic;
signal \n21948_cascade_\ : std_logic;
signal buf_adcdata_vac_22 : std_logic;
signal \AC_ADC_SYNC\ : std_logic;
signal \RTD.n21988\ : std_logic;
signal \RTD.n7_adj_1497_cascade_\ : std_logic;
signal \n13603_cascade_\ : std_logic;
signal read_buf_5 : std_logic;
signal \RTD.n62\ : std_logic;
signal \RTD.n12274\ : std_logic;
signal \RTD.n11_adj_1500\ : std_logic;
signal buf_adcdata_vac_23 : std_logic;
signal n23435 : std_logic;
signal \RTD.mode\ : std_logic;
signal \RTD.cfg_buf_6\ : std_logic;
signal \RTD.cfg_buf_5\ : std_logic;
signal \RTD.n12\ : std_logic;
signal \RTD.cfg_buf_1\ : std_logic;
signal \RTD.n20093\ : std_logic;
signal \RTD.n13482\ : std_logic;
signal \RTD.n68\ : std_logic;
signal \RTD.cfg_buf_7\ : std_logic;
signal \buf_readRTD_14\ : std_logic;
signal \RTD.n68_adj_1498\ : std_logic;
signal \RTD.n21954\ : std_logic;
signal \RTD_DRDY\ : std_logic;
signal \RTD.n21954_cascade_\ : std_logic;
signal \RTD.n21955\ : std_logic;
signal \RTD.adress_7_N_1009_7\ : std_logic;
signal \RTD.n11\ : std_logic;
signal \RTD.n11_cascade_\ : std_logic;
signal \RTD.n13488\ : std_logic;
signal \RTD.n13488_cascade_\ : std_logic;
signal \RTD.n15585\ : std_logic;
signal \RTD.n22081\ : std_logic;
signal \RTD.adress_6\ : std_logic;
signal \RTD.adress_5\ : std_logic;
signal \RTD.adress_4\ : std_logic;
signal \RTD.adress_3\ : std_logic;
signal \RTD.adress_2\ : std_logic;
signal \RTD.adress_0\ : std_logic;
signal \RTD.n13441\ : std_logic;
signal \RTD.adress_1\ : std_logic;
signal read_buf_6 : std_logic;
signal n21989 : std_logic;
signal n13584 : std_logic;
signal read_buf_7 : std_logic;
signal buf_adcdata_vac_9 : std_logic;
signal n19_adj_1752 : std_logic;
signal read_buf_8 : std_logic;
signal n13603 : std_logic;
signal read_buf_9 : std_logic;
signal \buf_readRTD_2\ : std_logic;
signal cmd_rdadctmp_12_adj_1536 : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal cmd_rdadctmp_22_adj_1526 : std_logic;
signal buf_adcdata_vac_15 : std_logic;
signal \n19_adj_1714_cascade_\ : std_logic;
signal \buf_readRTD_7\ : std_logic;
signal \CLK_DDS.tmp_buf_10\ : std_logic;
signal \CLK_DDS.tmp_buf_11\ : std_logic;
signal \CLK_DDS.tmp_buf_12\ : std_logic;
signal \CLK_DDS.tmp_buf_13\ : std_logic;
signal \CLK_DDS.tmp_buf_14\ : std_logic;
signal \CLK_DDS.tmp_buf_9\ : std_logic;
signal \CLK_DDS.tmp_buf_8\ : std_logic;
signal tmp_buf_15_adj_1511 : std_logic;
signal \CLK_DDS.tmp_buf_0\ : std_logic;
signal \CLK_DDS.tmp_buf_1\ : std_logic;
signal \CLK_DDS.tmp_buf_2\ : std_logic;
signal \CLK_DDS.tmp_buf_3\ : std_logic;
signal \CLK_DDS.tmp_buf_4\ : std_logic;
signal \CLK_DDS.tmp_buf_5\ : std_logic;
signal dds_state_2_adj_1508 : std_logic;
signal dds_state_1_adj_1509 : std_logic;
signal \CLK_DDS.tmp_buf_6\ : std_logic;
signal \CLK_DDS.tmp_buf_7\ : std_logic;
signal \CLK_DDS.n13376\ : std_logic;
signal n19_adj_1765 : std_logic;
signal n20_adj_1766 : std_logic;
signal \n21892_cascade_\ : std_logic;
signal \IAC_MISO\ : std_logic;
signal \GB_BUFFER_DDS_MCLK1_THRU_CO\ : std_logic;
signal n22388 : std_logic;
signal \VDC_SCLK\ : std_logic;
signal n12356 : std_logic;
signal \RTD.n17\ : std_logic;
signal \RTD.n79\ : std_logic;
signal buf_adcdata_vdc_15 : std_logic;
signal buf_adcdata_vdc_7 : std_logic;
signal buf_adcdata_vdc_23 : std_logic;
signal buf_adcdata_vdc_4 : std_logic;
signal buf_adcdata_vdc_9 : std_logic;
signal buf_adcdata_vdc_6 : std_logic;
signal buf_adcdata_vdc_22 : std_logic;
signal cmd_rdadctmp_26_adj_1522 : std_logic;
signal \n112_adj_1786_cascade_\ : std_logic;
signal buf_adcdata_vdc_10 : std_logic;
signal buf_adcdata_vac_10 : std_logic;
signal n19_adj_1747 : std_logic;
signal comm_test_buf_24_22 : std_logic;
signal buf_dds1_15 : std_logic;
signal n111_adj_1771 : std_logic;
signal buf_adcdata_vdc_8 : std_logic;
signal buf_adcdata_vac_8 : std_logic;
signal n30_adj_1695 : std_logic;
signal \buf_readRTD_11\ : std_logic;
signal \buf_cfgRTD_3\ : std_logic;
signal n20_adj_1790 : std_logic;
signal \n23498_cascade_\ : std_logic;
signal buf_adcdata_vdc_20 : std_logic;
signal buf_adcdata_vac_20 : std_logic;
signal n16_adj_1787 : std_logic;
signal n17_adj_1788 : std_logic;
signal n23540 : std_logic;
signal buf_adcdata_iac_23 : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal n19 : std_logic;
signal \buf_readRTD_0\ : std_logic;
signal \n22041_cascade_\ : std_logic;
signal \INVacadc_trig_303C_net\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \ADC_IAC.n20676\ : std_logic;
signal \ADC_IAC.n20677\ : std_logic;
signal \ADC_IAC.n20678\ : std_logic;
signal \ADC_IAC.n20679\ : std_logic;
signal \ADC_IAC.n20680\ : std_logic;
signal \ADC_IAC.n20681\ : std_logic;
signal \ADC_IAC.n20682\ : std_logic;
signal \ADC_IAC.n13667\ : std_logic;
signal \ADC_IAC.n15622\ : std_logic;
signal \ADC_IAC.n22031\ : std_logic;
signal \ADC_IAC.bit_cnt_4\ : std_logic;
signal \ADC_IAC.bit_cnt_3\ : std_logic;
signal \ADC_IAC.bit_cnt_1\ : std_logic;
signal \ADC_IAC.bit_cnt_2\ : std_logic;
signal \ADC_IAC.bit_cnt_6\ : std_logic;
signal \ADC_IAC.bit_cnt_0\ : std_logic;
signal \ADC_IAC.n22113_cascade_\ : std_logic;
signal \ADC_IAC.bit_cnt_7\ : std_logic;
signal \ADC_IAC.bit_cnt_5\ : std_logic;
signal \ADC_IAC.n22128_cascade_\ : std_logic;
signal \ADC_IAC.n22384_cascade_\ : std_logic;
signal \ADC_IAC.n22032\ : std_logic;
signal acadc_trig : std_logic;
signal \ADC_IAC.n17_cascade_\ : std_logic;
signal \ADC_IAC.n12\ : std_logic;
signal n21892 : std_logic;
signal n14_adj_1578 : std_logic;
signal \IAC_DRDY\ : std_logic;
signal \IAC_CS\ : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal \EIS_SYNCCLK\ : std_logic;
signal \IAC_CLK\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_1\ : std_logic;
signal \ADC_VDC.n20725\ : std_logic;
signal \ADC_VDC.avg_cnt_2\ : std_logic;
signal \ADC_VDC.n20726\ : std_logic;
signal \ADC_VDC.avg_cnt_3\ : std_logic;
signal \ADC_VDC.n20727\ : std_logic;
signal \ADC_VDC.avg_cnt_4\ : std_logic;
signal \ADC_VDC.n20728\ : std_logic;
signal \ADC_VDC.n20729\ : std_logic;
signal \ADC_VDC.avg_cnt_6\ : std_logic;
signal \ADC_VDC.n20730\ : std_logic;
signal \ADC_VDC.avg_cnt_7\ : std_logic;
signal \ADC_VDC.n20731\ : std_logic;
signal \ADC_VDC.n20732\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_9\ : std_logic;
signal \ADC_VDC.n20733\ : std_logic;
signal \ADC_VDC.n20734\ : std_logic;
signal \ADC_VDC.n20735\ : std_logic;
signal \ADC_VDC.avg_cnt_11\ : std_logic;
signal \RTD.adc_state_3\ : std_logic;
signal \RTD.adc_state_1\ : std_logic;
signal adc_state_2 : std_logic;
signal \RTD.adc_state_0\ : std_logic;
signal \ADC_VDC.n22071_cascade_\ : std_logic;
signal cmd_rdadctmp_0_adj_1574 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_0\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal cmd_rdadctmp_1_adj_1573 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_1\ : std_logic;
signal \ADC_VDC.n20690\ : std_logic;
signal cmd_rdadctmp_2_adj_1572 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_2\ : std_logic;
signal \ADC_VDC.n20691\ : std_logic;
signal cmd_rdadctmp_3_adj_1571 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_3\ : std_logic;
signal \ADC_VDC.n20692\ : std_logic;
signal cmd_rdadctmp_4_adj_1570 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_4\ : std_logic;
signal \ADC_VDC.n20693\ : std_logic;
signal cmd_rdadctmp_5_adj_1569 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_5\ : std_logic;
signal \ADC_VDC.n20694\ : std_logic;
signal cmd_rdadctmp_6_adj_1568 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_6\ : std_logic;
signal \ADC_VDC.n20695\ : std_logic;
signal cmd_rdadctmp_7_adj_1567 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_7\ : std_logic;
signal \ADC_VDC.n20696\ : std_logic;
signal \ADC_VDC.n20697\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_8\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_9\ : std_logic;
signal \ADC_VDC.n20698\ : std_logic;
signal cmd_rdadctmp_10_adj_1564 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_10\ : std_logic;
signal \ADC_VDC.n20699\ : std_logic;
signal cmd_rdadctmp_11_adj_1563 : std_logic;
signal \ADC_VDC.n20700\ : std_logic;
signal cmd_rdadctmp_12_adj_1562 : std_logic;
signal cmd_rdadcbuf_12 : std_logic;
signal \ADC_VDC.n20701\ : std_logic;
signal cmd_rdadctmp_13_adj_1561 : std_logic;
signal \ADC_VDC.n20702\ : std_logic;
signal cmd_rdadctmp_14_adj_1560 : std_logic;
signal \ADC_VDC.n20703\ : std_logic;
signal cmd_rdadctmp_15_adj_1559 : std_logic;
signal cmd_rdadcbuf_15 : std_logic;
signal \ADC_VDC.n20704\ : std_logic;
signal \ADC_VDC.n20705\ : std_logic;
signal cmd_rdadctmp_16_adj_1558 : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal cmd_rdadctmp_17_adj_1557 : std_logic;
signal cmd_rdadcbuf_17 : std_logic;
signal \ADC_VDC.n20706\ : std_logic;
signal cmd_rdadctmp_18_adj_1556 : std_logic;
signal cmd_rdadcbuf_18 : std_logic;
signal \ADC_VDC.n20707\ : std_logic;
signal cmd_rdadctmp_19_adj_1555 : std_logic;
signal cmd_rdadcbuf_19 : std_logic;
signal \ADC_VDC.n20708\ : std_logic;
signal cmd_rdadctmp_20_adj_1554 : std_logic;
signal cmd_rdadcbuf_20 : std_logic;
signal \ADC_VDC.n20709\ : std_logic;
signal cmd_rdadctmp_21_adj_1553 : std_logic;
signal cmd_rdadcbuf_21 : std_logic;
signal \ADC_VDC.n20710\ : std_logic;
signal \ADC_VDC.n20711\ : std_logic;
signal cmd_rdadcbuf_23 : std_logic;
signal \ADC_VDC.n20712\ : std_logic;
signal \ADC_VDC.n20713\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal cmd_rdadcbuf_25 : std_logic;
signal \ADC_VDC.n20714\ : std_logic;
signal cmd_rdadcbuf_26 : std_logic;
signal \ADC_VDC.n20715\ : std_logic;
signal \ADC_VDC.n20716\ : std_logic;
signal cmd_rdadcbuf_28 : std_logic;
signal \ADC_VDC.n20717\ : std_logic;
signal cmd_rdadcbuf_29 : std_logic;
signal \ADC_VDC.n20718\ : std_logic;
signal cmd_rdadcbuf_30 : std_logic;
signal \ADC_VDC.n20719\ : std_logic;
signal cmd_rdadcbuf_31 : std_logic;
signal \ADC_VDC.n20720\ : std_logic;
signal \ADC_VDC.n20721\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal cmd_rdadcbuf_33 : std_logic;
signal \ADC_VDC.n20722\ : std_logic;
signal \ADC_VDC.n20723\ : std_logic;
signal \n23474_cascade_\ : std_logic;
signal \n23477_cascade_\ : std_logic;
signal n30_adj_1784 : std_logic;
signal n112_adj_1772 : std_logic;
signal \n30_adj_1768_cascade_\ : std_logic;
signal n19_adj_1780 : std_logic;
signal n30_adj_1702 : std_logic;
signal n22358 : std_logic;
signal buf_adcdata_vdc_19 : std_logic;
signal n19_adj_1789 : std_logic;
signal n23426 : std_logic;
signal n23429 : std_logic;
signal cmd_rdadctmp_27_adj_1521 : std_logic;
signal buf_adcdata_vac_19 : std_logic;
signal buf_adcdata_iac_19 : std_logic;
signal buf_dds1_12 : std_logic;
signal n16_adj_1778 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal buf_dds1_7 : std_logic;
signal \IAC_SCLK\ : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal \ADC_VDC.avg_cnt_0\ : std_logic;
signal \ADC_VDC.avg_cnt_5\ : std_logic;
signal \ADC_VDC.avg_cnt_8\ : std_logic;
signal \ADC_VDC.avg_cnt_10\ : std_logic;
signal \ADC_VDC.n20\ : std_logic;
signal \ADC_VDC.n19_cascade_\ : std_logic;
signal \ADC_VDC.n21\ : std_logic;
signal \ADC_VDC.n28\ : std_logic;
signal \ADC_VDC.n21871\ : std_logic;
signal \ADC_VDC.n13865\ : std_logic;
signal \ADC_VDC.n9_cascade_\ : std_logic;
signal \ADC_VDC.n22071\ : std_logic;
signal \ADC_VDC.n5\ : std_logic;
signal cmd_rdadcbuf_14 : std_logic;
signal cmd_rdadctmp_8_adj_1566 : std_logic;
signal n13925 : std_logic;
signal cmd_rdadctmp_9_adj_1565 : std_logic;
signal cmd_rdadcbuf_22 : std_logic;
signal cmd_rdadcbuf_13 : std_logic;
signal cmd_rdadcbuf_16 : std_logic;
signal buf_adcdata_vdc_5 : std_logic;
signal cmd_rdadcbuf_27 : std_logic;
signal buf_dds1_5 : std_logic;
signal buf_adcdata_vdc_14 : std_logic;
signal buf_adcdata_vac_14 : std_logic;
signal \ADC_VDC.n14120\ : std_logic;
signal \ADC_VDC.n15721\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_35_N_1344_34\ : std_logic;
signal \ADC_VDC.n4_cascade_\ : std_logic;
signal cmd_rdadcbuf_34 : std_logic;
signal \ADC_VDC.n14092\ : std_logic;
signal \comm_spi.n24028\ : std_logic;
signal \comm_spi.n24028_cascade_\ : std_logic;
signal \buf_readRTD_12\ : std_logic;
signal n20_adj_1781 : std_logic;
signal cmd_rdadctmp_19_adj_1529 : std_logic;
signal cmd_rdadctmp_20_adj_1528 : std_logic;
signal n23309 : std_logic;
signal \buf_readRTD_10\ : std_logic;
signal \n22164_cascade_\ : std_logic;
signal buf_dds1_14 : std_logic;
signal n23366 : std_logic;
signal \n16_adj_1763_cascade_\ : std_logic;
signal n23369 : std_logic;
signal n30_adj_1698 : std_logic;
signal \buf_cfgRTD_6\ : std_logic;
signal \buf_cfgRTD_2\ : std_logic;
signal \buf_cfgRTD_4\ : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal buf_dds1_11 : std_logic;
signal data_count_0 : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n20613 : std_logic;
signal data_count_2 : std_logic;
signal n20614 : std_logic;
signal data_count_3 : std_logic;
signal n20615 : std_logic;
signal data_count_4 : std_logic;
signal n20616 : std_logic;
signal data_count_5 : std_logic;
signal n20617 : std_logic;
signal data_count_6 : std_logic;
signal n20618 : std_logic;
signal data_count_7 : std_logic;
signal n20619 : std_logic;
signal n20620 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal data_count_8 : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal n20621 : std_logic;
signal data_count_9 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal n11983 : std_logic;
signal \n24_adj_1598_cascade_\ : std_logic;
signal \n24_adj_1506_cascade_\ : std_logic;
signal \IAC_FLT1\ : std_logic;
signal n11982 : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal n23468 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal \DTRIG_N_1182\ : std_logic;
signal adc_state_1 : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal buf_adcdata_iac_17 : std_logic;
signal buf_dds1_10 : std_logic;
signal n22160 : std_logic;
signal buf_adcdata_iac_18 : std_logic;
signal \IAC_FLT0\ : std_logic;
signal n22161 : std_logic;
signal \ADC_VDC.adc_state_3_N_1316_1\ : std_logic;
signal \ADC_VDC.n22404_cascade_\ : std_logic;
signal \ADC_VDC.n17\ : std_logic;
signal \ADC_VDC.n17_cascade_\ : std_logic;
signal \ADC_VDC.n22055\ : std_logic;
signal \ADC_VDC.n27_cascade_\ : std_logic;
signal \ADC_VDC.n10\ : std_logic;
signal \ADC_VDC.n21869\ : std_logic;
signal \ADC_VDC.n11923\ : std_logic;
signal \ADC_VDC.n11923_cascade_\ : std_logic;
signal \ADC_VDC.n20869_cascade_\ : std_logic;
signal \ADC_VDC.n8031\ : std_logic;
signal \ADC_VDC.n23531\ : std_logic;
signal \ADC_VDC.n20869\ : std_logic;
signal \ADC_VDC.n21991\ : std_logic;
signal \ADC_VDC.n22075_cascade_\ : std_logic;
signal \ADC_VDC.n44_adj_1487\ : std_logic;
signal \ADC_VDC.n39_adj_1488\ : std_logic;
signal \ADC_VDC.n6_adj_1485\ : std_logic;
signal \ADC_VDC.n21859_cascade_\ : std_logic;
signal \ADC_VDC.n22628_cascade_\ : std_logic;
signal \ADC_VDC.n21859\ : std_logic;
signal \ADC_VDC.n22625\ : std_logic;
signal \ADC_VDC.n6\ : std_logic;
signal cmd_rdadctmp_22_adj_1552 : std_logic;
signal \ADC_VDC.n11183_cascade_\ : std_logic;
signal \ADC_VDC.cmd_rdadctmp_23\ : std_logic;
signal \ADC_VDC.n13957\ : std_logic;
signal \ADC_VDC.n21707\ : std_logic;
signal \INVcomm_spi.imiso_83_12612_12613_resetC_net\ : std_logic;
signal \comm_spi.n15369\ : std_logic;
signal \buf_readRTD_13\ : std_logic;
signal buf_adcdata_vac_21 : std_logic;
signal \buf_cfgRTD_5\ : std_logic;
signal \n23384_cascade_\ : std_logic;
signal cmd_rdadcbuf_32 : std_logic;
signal buf_adcdata_vdc_21 : std_logic;
signal cmd_rdadcbuf_24 : std_logic;
signal n12352 : std_logic;
signal cmd_rdadcbuf_11 : std_logic;
signal buf_adcdata_vdc_12 : std_logic;
signal buf_adcdata_vac_12 : std_logic;
signal \buf_readRTD_4\ : std_logic;
signal \n19_adj_1734_cascade_\ : std_logic;
signal cmd_rdadctmp_7_adj_1541 : std_logic;
signal cmd_rdadctmp_6_adj_1542 : std_logic;
signal cmd_rdadctmp_5_adj_1543 : std_logic;
signal cmd_rdadctmp_3_adj_1545 : std_logic;
signal cmd_rdadctmp_4_adj_1544 : std_logic;
signal buf_dds1_6 : std_logic;
signal buf_data_iac_0 : std_logic;
signal cmd_rdadctmp_21_adj_1527 : std_logic;
signal n30_adj_1692 : std_logic;
signal cmd_rdadctmp_25_adj_1523 : std_logic;
signal buf_adcdata_vdc_18 : std_logic;
signal buf_adcdata_vac_18 : std_logic;
signal n22163 : std_logic;
signal \comm_spi.n15360\ : std_logic;
signal \comm_spi.data_tx_7__N_857\ : std_logic;
signal comm_test_buf_24_19 : std_logic;
signal comm_test_buf_24_20 : std_logic;
signal n111_adj_1785 : std_logic;
signal \n24_cascade_\ : std_logic;
signal buf_adcdata_iac_22 : std_logic;
signal \VAC_FLT0\ : std_logic;
signal n17_adj_1764 : std_logic;
signal \n11981_cascade_\ : std_logic;
signal \VAC_FLT1\ : std_logic;
signal n24_adj_1576 : std_logic;
signal n11986 : std_logic;
signal \n23510_cascade_\ : std_logic;
signal n22276 : std_logic;
signal \n23513_cascade_\ : std_logic;
signal \n30_adj_1759_cascade_\ : std_logic;
signal n26_adj_1758 : std_logic;
signal eis_end : std_logic;
signal \INVeis_end_302C_net\ : std_logic;
signal n112_adj_1762 : std_logic;
signal \n21946_cascade_\ : std_logic;
signal n21880 : std_logic;
signal \n13_cascade_\ : std_logic;
signal \INVeis_state_i2C_net\ : std_logic;
signal n22395 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal n13_adj_1591 : std_logic;
signal n11_adj_1592 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal acadc_dtrig_i : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal \DTRIG_N_1182_adj_1549\ : std_logic;
signal adc_state_1_adj_1515 : std_logic;
signal acadc_dtrig_v : std_logic;
signal buf_dds1_9 : std_logic;
signal n23534 : std_logic;
signal buf_dds0_10 : std_logic;
signal buf_dds0_6 : std_logic;
signal buf_dds0_5 : std_logic;
signal \SIG_DDS.tmp_buf_4\ : std_logic;
signal \SIG_DDS.tmp_buf_5\ : std_logic;
signal \SIG_DDS.tmp_buf_9\ : std_logic;
signal \SIG_DDS.tmp_buf_6\ : std_logic;
signal buf_dds0_7 : std_logic;
signal buf_dds0_12 : std_logic;
signal \SIG_DDS.tmp_buf_12\ : std_logic;
signal \SIG_DDS.tmp_buf_13\ : std_logic;
signal buf_dds0_14 : std_logic;
signal \SIG_DDS.tmp_buf_14\ : std_logic;
signal buf_dds0_15 : std_logic;
signal \SIG_DDS.tmp_buf_7\ : std_logic;
signal \SIG_DDS.tmp_buf_8\ : std_logic;
signal \SIG_DDS.tmp_buf_10\ : std_logic;
signal buf_dds0_11 : std_logic;
signal \SIG_DDS.tmp_buf_11\ : std_logic;
signal \ADC_VDC.n22063\ : std_logic;
signal \RTD.n20050\ : std_logic;
signal \VDC_SDO\ : std_logic;
signal \ADC_VDC.n35_cascade_\ : std_logic;
signal \ADC_VDC.n45\ : std_logic;
signal \ADC_VDC.n22067\ : std_logic;
signal adc_state_3 : std_logic;
signal adc_state_1_adj_1551 : std_logic;
signal \ADC_VDC.adc_state_0\ : std_logic;
signal adc_state_2_adj_1550 : std_logic;
signal \ADC_VDC.n11183\ : std_logic;
signal \ADC_VDC.n23528\ : std_logic;
signal \ADC_VDC.bit_cnt_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \ADC_VDC.bit_cnt_1\ : std_logic;
signal \ADC_VDC.n20812\ : std_logic;
signal \ADC_VDC.bit_cnt_2\ : std_logic;
signal \ADC_VDC.n20813\ : std_logic;
signal \ADC_VDC.bit_cnt_3\ : std_logic;
signal \ADC_VDC.n20814\ : std_logic;
signal \ADC_VDC.bit_cnt_4\ : std_logic;
signal \ADC_VDC.n20815\ : std_logic;
signal \ADC_VDC.bit_cnt_5\ : std_logic;
signal \ADC_VDC.n20816\ : std_logic;
signal \ADC_VDC.bit_cnt_6\ : std_logic;
signal \ADC_VDC.n20817\ : std_logic;
signal \ADC_VDC.n20818\ : std_logic;
signal \ADC_VDC.bit_cnt_7\ : std_logic;
signal \ADC_VDC.n17565\ : std_logic;
signal \ADC_VDC.n17542\ : std_logic;
signal \comm_spi.n15361\ : std_logic;
signal buf_adcdata_vdc_3 : std_logic;
signal \n19_adj_1703_cascade_\ : std_logic;
signal buf_data_iac_3 : std_logic;
signal \n22_adj_1704_cascade_\ : std_logic;
signal buf_adcdata_iac_3 : std_logic;
signal cmd_rdadctmp_11_adj_1537 : std_logic;
signal buf_adcdata_vac_3 : std_logic;
signal buf_adcdata_vdc_1 : std_logic;
signal buf_adcdata_vac_1 : std_logic;
signal \n19_adj_1710_cascade_\ : std_logic;
signal buf_data_iac_1 : std_logic;
signal \n22_adj_1711_cascade_\ : std_logic;
signal \n30_adj_1712_cascade_\ : std_logic;
signal \comm_spi.n24031\ : std_logic;
signal n30_adj_1705 : std_logic;
signal n13847 : std_logic;
signal cmd_rdadctmp_9_adj_1539 : std_logic;
signal \n2_adj_1666_cascade_\ : std_logic;
signal n1_adj_1665 : std_logic;
signal \comm_spi.data_tx_7__N_865\ : std_logic;
signal comm_test_buf_24_4 : std_logic;
signal n13231 : std_logic;
signal n13237 : std_logic;
signal n22295 : std_logic;
signal n4_adj_1667 : std_logic;
signal n23294 : std_logic;
signal n30_adj_1588 : std_logic;
signal comm_test_buf_24_3 : std_logic;
signal n111_adj_1794 : std_logic;
signal n15545 : std_logic;
signal buf_dds1_8 : std_logic;
signal comm_test_buf_24_11 : std_logic;
signal comm_test_buf_24_12 : std_logic;
signal buf_adcdata_iac_16 : std_logic;
signal n23324 : std_logic;
signal req_data_cnt_8 : std_logic;
signal \n19_adj_1727_cascade_\ : std_logic;
signal \n29_adj_1770_cascade_\ : std_logic;
signal comm_test_buf_24_14 : std_logic;
signal comm_test_buf_24_6 : std_logic;
signal n16_adj_1683 : std_logic;
signal \n17642_cascade_\ : std_logic;
signal n22312 : std_logic;
signal n23330 : std_logic;
signal n17633 : std_logic;
signal \iac_raw_buf_N_821\ : std_logic;
signal n17_adj_1742 : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal n12369 : std_logic;
signal n24_adj_1503 : std_logic;
signal n11980 : std_logic;
signal eis_state_0 : std_logic;
signal eis_state_2 : std_logic;
signal \n12450_cascade_\ : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n22120 : std_logic;
signal n20637 : std_logic;
signal \n20637_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n20637_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n20637_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n20637_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n20637_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n20637_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n20637_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal n20638 : std_logic;
signal n20639 : std_logic;
signal n20640 : std_logic;
signal n20641 : std_logic;
signal n20642 : std_logic;
signal n20643 : std_logic;
signal n20644 : std_logic;
signal n20645 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal n20646 : std_logic;
signal n20647 : std_logic;
signal n20648 : std_logic;
signal n20649 : std_logic;
signal n20650 : std_logic;
signal n20651 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal n12450 : std_logic;
signal n15439 : std_logic;
signal \RTD.bit_cnt_3\ : std_logic;
signal \RTD.bit_cnt_2\ : std_logic;
signal \RTD.bit_cnt_1\ : std_logic;
signal \RTD.bit_cnt_0\ : std_logic;
signal \clk_RTD\ : std_logic;
signal \RTD.n18274\ : std_logic;
signal \RTD.n18275\ : std_logic;
signal \buf_cfgRTD_7\ : std_logic;
signal \buf_readRTD_15\ : std_logic;
signal n23432 : std_logic;
signal \n12610_cascade_\ : std_logic;
signal \comm_spi.data_tx_7__N_883\ : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \comm_spi.data_tx_7__N_868\ : std_logic;
signal buf_adcdata_vdc_2 : std_logic;
signal \n19_adj_1706_cascade_\ : std_logic;
signal cmd_rdadctmp_8_adj_1540 : std_logic;
signal buf_adcdata_iac_1 : std_logic;
signal buf_adcdata_iac_2 : std_logic;
signal cmd_rdadctmp_10_adj_1538 : std_logic;
signal adc_state_0_adj_1516 : std_logic;
signal n21948 : std_logic;
signal buf_adcdata_vac_2 : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal \comm_spi.n24034_cascade_\ : std_logic;
signal \comm_spi.n15356\ : std_logic;
signal \comm_spi.data_tx_7__N_858\ : std_logic;
signal comm_tx_buf_6 : std_logic;
signal \comm_spi.n24013\ : std_logic;
signal \comm_spi.data_tx_7__N_856\ : std_logic;
signal \n2_adj_1669_cascade_\ : std_logic;
signal \n4_adj_1670_cascade_\ : std_logic;
signal n23402 : std_logic;
signal n22669 : std_logic;
signal n1_adj_1668 : std_logic;
signal n13219 : std_logic;
signal comm_tx_buf_4 : std_logic;
signal \comm_spi.data_tx_7__N_871\ : std_logic;
signal \comm_buf_0_7_N_543_4\ : std_logic;
signal \comm_buf_0_7_N_543_6\ : std_logic;
signal \comm_buf_0_7_N_543_7\ : std_logic;
signal clk_cnt_1 : std_logic;
signal clk_cnt_0 : std_logic;
signal n18996 : std_logic;
signal \comm_buf_2_7_N_575_0\ : std_logic;
signal \comm_buf_2_7_N_575_1\ : std_logic;
signal \comm_buf_2_7_N_575_3\ : std_logic;
signal \comm_buf_2_7_N_575_4\ : std_logic;
signal \comm_buf_2_7_N_575_5\ : std_logic;
signal \comm_buf_2_7_N_575_6\ : std_logic;
signal comm_buf_2_6 : std_logic;
signal \comm_buf_2_7_N_575_7\ : std_logic;
signal \comm_spi.data_tx_7__N_859\ : std_logic;
signal n6774 : std_logic;
signal \n111_adj_1796_cascade_\ : std_logic;
signal comm_test_buf_24_10 : std_logic;
signal \comm_spi.n15365\ : std_logic;
signal \comm_spi.n24025\ : std_logic;
signal \comm_spi.n15364\ : std_logic;
signal \comm_spi.n15368\ : std_logic;
signal \comm_spi.data_tx_7__N_855\ : std_logic;
signal \AMPV_POW\ : std_logic;
signal n111_adj_1761 : std_logic;
signal buf_dds1_3 : std_logic;
signal comm_buf_2_4 : std_logic;
signal \n11987_cascade_\ : std_logic;
signal n17_adj_1779 : std_logic;
signal \n11985_cascade_\ : std_logic;
signal n13117 : std_logic;
signal n15538 : std_logic;
signal \IAC_OSR0\ : std_logic;
signal n24_adj_1575 : std_logic;
signal \IAC_OSR1\ : std_logic;
signal n24_adj_1601 : std_logic;
signal n11984 : std_logic;
signal n16_adj_1733 : std_logic;
signal n23438 : std_logic;
signal buf_adcdata_iac_12 : std_logic;
signal comm_test_buf_24_21 : std_logic;
signal comm_test_buf_24_13 : std_logic;
signal comm_test_buf_24_5 : std_logic;
signal \n111_adj_1776_cascade_\ : std_logic;
signal n11979 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal buf_dds1_0 : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal buf_adcdata_iac_20 : std_logic;
signal buf_control_6 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal n23_adj_1767 : std_logic;
signal \SIG_DDS.tmp_buf_0\ : std_logic;
signal \SIG_DDS.tmp_buf_3\ : std_logic;
signal \SIG_DDS.tmp_buf_1\ : std_logic;
signal \SIG_DDS.tmp_buf_2\ : std_logic;
signal \comm_spi.n15323\ : std_logic;
signal \comm_spi.data_tx_7__N_860\ : std_logic;
signal \comm_spi.n24040\ : std_logic;
signal \comm_spi.data_tx_7__N_880\ : std_logic;
signal \comm_spi.n24037\ : std_logic;
signal \comm_spi.n15348\ : std_logic;
signal \comm_spi.n15349\ : std_logic;
signal \comm_spi.n15335\ : std_logic;
signal \INVcomm_spi.MISO_48_12606_12607_resetC_net\ : std_logic;
signal n23390 : std_logic;
signal \n1_adj_1674_cascade_\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal n22341 : std_logic;
signal n2_adj_1675 : std_logic;
signal buf_adcdata_vdc_0 : std_logic;
signal buf_adcdata_vac_0 : std_logic;
signal \n19_adj_1590_cascade_\ : std_logic;
signal n22_adj_1589 : std_logic;
signal \n21965_cascade_\ : std_logic;
signal n13746 : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal comm_buf_6_4 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal buf_adcdata_iac_0 : std_logic;
signal buf_adcdata_vdc_13 : std_logic;
signal buf_adcdata_vac_13 : std_logic;
signal \buf_readRTD_5\ : std_logic;
signal \n19_adj_1729_cascade_\ : std_logic;
signal comm_buf_6_6 : std_logic;
signal \n9_adj_1600_cascade_\ : std_logic;
signal \n6776_cascade_\ : std_logic;
signal n18890 : std_logic;
signal comm_test_buf_24_9 : std_logic;
signal \comm_buf_0_7_N_543_0\ : std_logic;
signal comm_test_buf_24_18 : std_logic;
signal comm_test_buf_24_7 : std_logic;
signal comm_test_buf_24_15 : std_logic;
signal comm_buf_2_1 : std_logic;
signal n13201 : std_logic;
signal \buf_readRTD_9\ : std_logic;
signal \buf_cfgRTD_1\ : std_logic;
signal \comm_spi.n15337\ : std_logic;
signal \comm_spi.n15338\ : std_logic;
signal \INVcomm_spi.imiso_83_12612_12613_setC_net\ : std_logic;
signal n15496 : std_logic;
signal buf_data_iac_16 : std_logic;
signal \n22270_cascade_\ : std_logic;
signal \n23450_cascade_\ : std_logic;
signal n23327 : std_logic;
signal n23453 : std_logic;
signal n112_adj_1583 : std_logic;
signal n23522 : std_logic;
signal n22267 : std_logic;
signal n112_adj_1797 : std_logic;
signal \comm_buf_0_7_N_543_2\ : std_logic;
signal comm_test_buf_24_16 : std_logic;
signal n111_adj_1584 : std_logic;
signal n20_adj_1804 : std_logic;
signal req_data_cnt_12 : std_logic;
signal \VAC_OSR1\ : std_logic;
signal buf_adcdata_iac_21 : std_logic;
signal n9_adj_1600 : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal n20652 : std_logic;
signal n20653 : std_logic;
signal n20654 : std_logic;
signal n20655 : std_logic;
signal n20656 : std_logic;
signal n20657 : std_logic;
signal n20658 : std_logic;
signal n20659 : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal n20660 : std_logic;
signal eis_stop : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal \VAC_OSR0\ : std_logic;
signal n40 : std_logic;
signal n24_adj_1505 : std_logic;
signal req_data_cnt_10 : std_logic;
signal acadc_rst : std_logic;
signal \data_index_9_N_236_3\ : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal n23_adj_1514 : std_logic;
signal n24_adj_1513 : std_logic;
signal \n21_cascade_\ : std_logic;
signal n22 : std_logic;
signal \n14_adj_1610_cascade_\ : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal \SELIRNG0\ : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal \VDC_RNG0\ : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal n23_adj_1783 : std_logic;
signal adc_state_0 : std_logic;
signal n21951 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal buf_dds0_8 : std_logic;
signal data_index_1 : std_logic;
signal n8_adj_1630 : std_logic;
signal \n8_adj_1630_cascade_\ : std_logic;
signal n7_adj_1629 : std_logic;
signal \data_index_9_N_236_1\ : std_logic;
signal buf_dds0_3 : std_logic;
signal tmp_buf_15 : std_logic;
signal \DDS_MOSI\ : std_logic;
signal \comm_spi.n24016\ : std_logic;
signal \comm_spi.n15326\ : std_logic;
signal \comm_spi.n24016_cascade_\ : std_logic;
signal \comm_spi.n15322\ : std_logic;
signal \comm_spi.data_tx_7__N_861\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal n20790 : std_logic;
signal n20791 : std_logic;
signal n20792 : std_logic;
signal n20793 : std_logic;
signal n20794 : std_logic;
signal n20795 : std_logic;
signal n20796 : std_logic;
signal n20797 : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal n20798 : std_logic;
signal n20799 : std_logic;
signal n20800 : std_logic;
signal n20801 : std_logic;
signal n20802 : std_logic;
signal n20803 : std_logic;
signal n20804 : std_logic;
signal n20805 : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal n20806 : std_logic;
signal n20807 : std_logic;
signal n20808 : std_logic;
signal n20809 : std_logic;
signal n20810 : std_logic;
signal n20811 : std_logic;
signal secclk_cnt_19 : std_logic;
signal secclk_cnt_21 : std_logic;
signal secclk_cnt_12 : std_logic;
signal secclk_cnt_22 : std_logic;
signal comm_buf_0_6 : std_logic;
signal comm_buf_6_1 : std_logic;
signal buf_data_iac_2 : std_logic;
signal n22_adj_1707 : std_logic;
signal comm_buf_2_7 : std_logic;
signal \n22331_cascade_\ : std_logic;
signal \n23360_cascade_\ : std_logic;
signal n2_adj_1663 : std_logic;
signal n4_adj_1664 : std_logic;
signal n1 : std_logic;
signal comm_tx_buf_7 : std_logic;
signal \comm_spi.data_tx_7__N_862\ : std_logic;
signal n4_adj_1673 : std_logic;
signal \n22342_cascade_\ : std_logic;
signal n23396 : std_logic;
signal \n1_adj_1671_cascade_\ : std_logic;
signal n2_adj_1672 : std_logic;
signal comm_buf_2_2 : std_logic;
signal comm_buf_0_2 : std_logic;
signal n13207 : std_logic;
signal comm_tx_buf_2 : std_logic;
signal \comm_spi.data_tx_7__N_877\ : std_logic;
signal buf_data_vac_16 : std_logic;
signal buf_data_vac_23 : std_logic;
signal comm_buf_3_7 : std_logic;
signal buf_data_vac_22 : std_logic;
signal comm_buf_3_6 : std_logic;
signal buf_data_vac_21 : std_logic;
signal buf_data_vac_20 : std_logic;
signal comm_buf_3_4 : std_logic;
signal buf_data_vac_19 : std_logic;
signal buf_data_vac_18 : std_logic;
signal comm_buf_3_2 : std_logic;
signal buf_data_vac_17 : std_logic;
signal comm_buf_3_1 : std_logic;
signal n15503 : std_logic;
signal n30_adj_1708 : std_logic;
signal comm_test_buf_24_2 : std_logic;
signal \comm_buf_2_7_N_575_2\ : std_logic;
signal n12880 : std_logic;
signal n21886 : std_logic;
signal \n12_cascade_\ : std_logic;
signal n15553 : std_logic;
signal n16_adj_1721 : std_logic;
signal buf_adcdata_iac_14 : std_logic;
signal n12015 : std_logic;
signal \n8_cascade_\ : std_logic;
signal buf_adcdata_vdc_11 : std_logic;
signal buf_adcdata_vac_11 : std_logic;
signal n22092 : std_logic;
signal n13211 : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal n23_adj_1756 : std_logic;
signal n21_adj_1803 : std_logic;
signal n30_adj_1769 : std_logic;
signal n22167 : std_logic;
signal n22166 : std_logic;
signal n23471 : std_logic;
signal \n23549_cascade_\ : std_logic;
signal n22174 : std_logic;
signal n112 : std_logic;
signal n30_adj_1805 : std_logic;
signal n17650 : std_logic;
signal n12 : std_logic;
signal buf_data_iac_12 : std_logic;
signal data_index_2 : std_logic;
signal n8_adj_1628 : std_logic;
signal \n8_adj_1628_cascade_\ : std_logic;
signal n7_adj_1627 : std_logic;
signal \data_index_9_N_236_2\ : std_logic;
signal n18865 : std_logic;
signal n7_adj_1626 : std_logic;
signal data_index_3 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal n20 : std_logic;
signal n14_adj_1599 : std_logic;
signal n17 : std_logic;
signal \n26_cascade_\ : std_logic;
signal n30_adj_1743 : std_logic;
signal n31 : std_logic;
signal buf_dds0_1 : std_logic;
signal buf_dds1_1 : std_logic;
signal buf_dds1_2 : std_logic;
signal buf_adcdata_iac_10 : std_logic;
signal \n16_adj_1746_cascade_\ : std_logic;
signal \comm_spi.n15341\ : std_logic;
signal \comm_spi.n15340\ : std_logic;
signal \comm_spi.n15333\ : std_logic;
signal \comm_spi.n15334\ : std_logic;
signal \INVcomm_spi.MISO_48_12606_12607_setC_net\ : std_logic;
signal \comm_spi.data_tx_7__N_854\ : std_logic;
signal comm_test_buf_24_1 : std_logic;
signal n111_adj_1798 : std_logic;
signal n21965 : std_logic;
signal \n12056_cascade_\ : std_logic;
signal comm_test_buf_24_23 : std_logic;
signal buf_dds0_2 : std_logic;
signal data_index_9 : std_logic;
signal \n8_adj_1617_cascade_\ : std_logic;
signal \data_index_9_N_236_8\ : std_logic;
signal \SIG_DDS.n13338\ : std_logic;
signal \comm_spi.iclk_N_850\ : std_logic;
signal \comm_spi.n15327\ : std_logic;
signal \VDC_CLK\ : std_logic;
signal \INVADC_VDC.genclk.t_clk_24C_net\ : std_logic;
signal n4_adj_1676 : std_logic;
signal \comm_spi.DOUT_7__N_835\ : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.iclk_N_851\ : std_logic;
signal secclk_cnt_15 : std_logic;
signal secclk_cnt_8 : std_logic;
signal secclk_cnt_1 : std_logic;
signal secclk_cnt_5 : std_logic;
signal \n25_adj_1717_cascade_\ : std_logic;
signal secclk_cnt_20 : std_logic;
signal \n20922_cascade_\ : std_logic;
signal n14_adj_1678 : std_logic;
signal secclk_cnt_9 : std_logic;
signal secclk_cnt_17 : std_logic;
signal n10_adj_1679 : std_logic;
signal secclk_cnt_6 : std_logic;
signal secclk_cnt_14 : std_logic;
signal secclk_cnt_10 : std_logic;
signal secclk_cnt_3 : std_logic;
signal n27 : std_logic;
signal secclk_cnt_16 : std_logic;
signal secclk_cnt_7 : std_logic;
signal secclk_cnt_13 : std_logic;
signal secclk_cnt_2 : std_logic;
signal n26_adj_1715 : std_logic;
signal n15420 : std_logic;
signal \TEST_LED\ : std_logic;
signal n9_adj_1596 : std_logic;
signal comm_buf_6_7 : std_logic;
signal comm_test_buf_24_17 : std_logic;
signal comm_buf_6_0 : std_logic;
signal \n18818_cascade_\ : std_logic;
signal \n23372_cascade_\ : std_logic;
signal n18816 : std_logic;
signal comm_tx_buf_0 : std_logic;
signal comm_buf_3_0 : std_logic;
signal n22338 : std_logic;
signal n18815 : std_logic;
signal comm_buf_2_0 : std_logic;
signal n18823 : std_logic;
signal buf_data_vac_0 : std_logic;
signal comm_buf_5_0 : std_logic;
signal buf_data_vac_7 : std_logic;
signal comm_buf_5_7 : std_logic;
signal buf_data_vac_6 : std_logic;
signal comm_buf_5_6 : std_logic;
signal buf_data_vac_5 : std_logic;
signal buf_data_vac_4 : std_logic;
signal comm_buf_5_4 : std_logic;
signal buf_data_vac_3 : std_logic;
signal buf_data_vac_2 : std_logic;
signal comm_buf_5_2 : std_logic;
signal buf_data_vac_1 : std_logic;
signal comm_buf_5_1 : std_logic;
signal \buf_readRTD_8\ : std_logic;
signal buf_adcdata_vdc_16 : std_logic;
signal \n23504_cascade_\ : std_logic;
signal buf_adcdata_vac_16 : std_logic;
signal n22288 : std_logic;
signal n12838 : std_logic;
signal n23306 : std_logic;
signal n8_adj_1504 : std_logic;
signal \n6_cascade_\ : std_logic;
signal n21938 : std_logic;
signal n19_adj_1722 : std_logic;
signal \buf_readRTD_6\ : std_logic;
signal n23288 : std_logic;
signal \n22396_cascade_\ : std_logic;
signal n6 : std_logic;
signal n22061 : std_logic;
signal n21929 : std_logic;
signal n22_adj_1801 : std_logic;
signal n112_adj_1799 : std_logic;
signal \comm_buf_0_7_N_543_1\ : std_logic;
signal n18_adj_1699 : std_logic;
signal n13257 : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n18 : std_logic;
signal comm_buf_0_0 : std_logic;
signal n11172 : std_logic;
signal eis_start : std_logic;
signal \n8_adj_1625_cascade_\ : std_logic;
signal \data_index_9_N_236_4\ : std_logic;
signal n7_adj_1624 : std_logic;
signal n8_adj_1625 : std_logic;
signal data_index_4 : std_logic;
signal n23546 : std_logic;
signal n30 : std_logic;
signal n17_adj_1594 : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal n24_adj_1800 : std_logic;
signal req_data_cnt_9 : std_logic;
signal req_data_cnt_15 : std_logic;
signal n22314 : std_logic;
signal n22169 : std_logic;
signal req_data_cnt_3 : std_logic;
signal \n23312_cascade_\ : std_logic;
signal \n23315_cascade_\ : std_logic;
signal n111_adj_1744 : std_logic;
signal \n30_adj_1741_cascade_\ : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal n19_adj_1739 : std_logic;
signal \buf_readRTD_3\ : std_logic;
signal buf_adcdata_iac_11 : std_logic;
signal n16_adj_1738 : std_logic;
signal \n23558_cascade_\ : std_logic;
signal n23561 : std_logic;
signal \SIG_DDS.bit_cnt_2\ : std_logic;
signal \SIG_DDS.bit_cnt_1\ : std_logic;
signal comm_buf_0_4 : std_logic;
signal comm_buf_0_1 : std_logic;
signal \SIG_DDS.bit_cnt_3\ : std_logic;
signal n8_adj_1615 : std_logic;
signal n7_adj_1614 : std_logic;
signal \data_index_9_N_236_9\ : std_logic;
signal data_index_6 : std_logic;
signal n8_adj_1621 : std_logic;
signal \n8_adj_1621_cascade_\ : std_logic;
signal n7_adj_1620 : std_logic;
signal \data_index_9_N_236_6\ : std_logic;
signal data_index_7 : std_logic;
signal n8_adj_1617 : std_logic;
signal n7_adj_1616 : std_logic;
signal data_index_8 : std_logic;
signal n8_adj_1619 : std_logic;
signal n7_adj_1618 : std_logic;
signal \data_index_9_N_236_7\ : std_logic;
signal \SIG_DDS.n22671\ : std_logic;
signal \SIG_DDS.n10\ : std_logic;
signal \comm_spi.imosi_N_841\ : std_logic;
signal \comm_spi.n15331\ : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.n24019\ : std_logic;
signal \comm_spi.n15344\ : std_logic;
signal \comm_spi.n15345\ : std_logic;
signal \comm_spi.n24019_cascade_\ : std_logic;
signal secclk_cnt_0 : std_logic;
signal secclk_cnt_18 : std_logic;
signal secclk_cnt_11 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n28 : std_logic;
signal \n12_adj_1760_cascade_\ : std_logic;
signal \n20834_cascade_\ : std_logic;
signal n30_adj_1681 : std_logic;
signal n33 : std_logic;
signal n32 : std_logic;
signal \n34_cascade_\ : std_logic;
signal n31_adj_1680 : std_logic;
signal \n49_cascade_\ : std_logic;
signal \comm_spi.n24022\ : std_logic;
signal \n8856_cascade_\ : std_logic;
signal n13273 : std_logic;
signal comm_buf_0_5 : std_logic;
signal comm_buf_3_5 : std_logic;
signal comm_buf_6_5 : std_logic;
signal comm_buf_2_5 : std_logic;
signal n18882 : std_logic;
signal \n18883_cascade_\ : std_logic;
signal comm_tx_buf_5 : std_logic;
signal comm_buf_5_5 : std_logic;
signal n22371 : std_logic;
signal \n18885_cascade_\ : std_logic;
signal n23414 : std_logic;
signal n22618 : std_logic;
signal n8_adj_1755 : std_logic;
signal n12976 : std_logic;
signal \n12976_cascade_\ : std_logic;
signal comm_buf_6_2 : std_logic;
signal \n22375_cascade_\ : std_logic;
signal buf_data_iac_22 : std_logic;
signal n22297 : std_logic;
signal \INVcomm_spi.bit_cnt_3787__i3C_net\ : std_logic;
signal eis_state_1 : std_logic;
signal n15517 : std_logic;
signal n12585 : std_logic;
signal n15238 : std_logic;
signal n12958 : std_logic;
signal n22397 : std_logic;
signal n29_adj_1688 : std_logic;
signal \n11402_cascade_\ : std_logic;
signal \comm_state_3_N_500_2\ : std_logic;
signal \n18850_cascade_\ : std_logic;
signal n13076 : std_logic;
signal n15531 : std_logic;
signal comm_buf_3_3 : std_logic;
signal comm_buf_6_3 : std_logic;
signal n18851 : std_logic;
signal comm_buf_5_3 : std_logic;
signal n22346 : std_logic;
signal \n18853_cascade_\ : std_logic;
signal n23378 : std_logic;
signal n6776 : std_logic;
signal comm_buf_2_3 : std_logic;
signal n18858 : std_logic;
signal comm_tx_buf_3 : std_logic;
signal \THERMOSTAT\ : std_logic;
signal buf_control_7 : std_logic;
signal \n12021_cascade_\ : std_logic;
signal n12614 : std_logic;
signal \n25_cascade_\ : std_logic;
signal n12548 : std_logic;
signal comm_buf_0_7 : std_logic;
signal n21964 : std_logic;
signal n11379 : std_logic;
signal n9 : std_logic;
signal n22059 : std_logic;
signal n26_adj_1740 : std_logic;
signal \n26_adj_1580_cascade_\ : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal \n23552_cascade_\ : std_logic;
signal req_data_cnt_0 : std_logic;
signal n16 : std_logic;
signal n23300 : std_logic;
signal buf_adcdata_iac_8 : std_logic;
signal buf_adcdata_iac_15 : std_logic;
signal n16_adj_1713 : std_logic;
signal n22268 : std_logic;
signal n13141 : std_logic;
signal n12610 : std_logic;
signal buf_dds0_4 : std_logic;
signal buf_dds0_0 : std_logic;
signal data_idxvec_0 : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal n14_adj_1613 : std_logic;
signal n20661 : std_logic;
signal n14_adj_1612 : std_logic;
signal n20662 : std_logic;
signal data_idxvec_3 : std_logic;
signal n20663 : std_logic;
signal n20664 : std_logic;
signal n14_adj_1661 : std_logic;
signal n20665 : std_logic;
signal n14_adj_1610 : std_logic;
signal n20666 : std_logic;
signal n14_adj_1609 : std_logic;
signal n20667 : std_logic;
signal n20668 : std_logic;
signal data_idxvec_8 : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal n20669 : std_logic;
signal n14_adj_1655 : std_logic;
signal data_idxvec_10 : std_logic;
signal n20670 : std_logic;
signal n20671 : std_logic;
signal n14_adj_1653 : std_logic;
signal n20672 : std_logic;
signal n20673 : std_logic;
signal n20674 : std_logic;
signal n14_adj_1607 : std_logic;
signal n20675 : std_logic;
signal data_idxvec_15 : std_logic;
signal data_index_0 : std_logic;
signal n11254 : std_logic;
signal n13052 : std_logic;
signal n15562 : std_logic;
signal \n15562_cascade_\ : std_logic;
signal bit_cnt_0 : std_logic;
signal \SIG_DDS.n9\ : std_logic;
signal \DDS_SCK\ : std_logic;
signal trig_dds0 : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.DOUT_7__N_834\ : std_logic;
signal \comm_spi.n15330\ : std_logic;
signal wdtick_cnt_0 : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal wdtick_cnt_1 : std_logic;
signal n20766 : std_logic;
signal wdtick_cnt_2 : std_logic;
signal n20767 : std_logic;
signal wdtick_cnt_3 : std_logic;
signal n20768 : std_logic;
signal wdtick_cnt_4 : std_logic;
signal n20769 : std_logic;
signal wdtick_cnt_5 : std_logic;
signal n20770 : std_logic;
signal wdtick_cnt_6 : std_logic;
signal n20771 : std_logic;
signal wdtick_cnt_7 : std_logic;
signal n20772 : std_logic;
signal n20773 : std_logic;
signal wdtick_cnt_8 : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal wdtick_cnt_9 : std_logic;
signal n20774 : std_logic;
signal wdtick_cnt_10 : std_logic;
signal n20775 : std_logic;
signal wdtick_cnt_11 : std_logic;
signal n20776 : std_logic;
signal wdtick_cnt_12 : std_logic;
signal n20777 : std_logic;
signal wdtick_cnt_13 : std_logic;
signal n20778 : std_logic;
signal wdtick_cnt_14 : std_logic;
signal n20779 : std_logic;
signal wdtick_cnt_15 : std_logic;
signal n20780 : std_logic;
signal n20781 : std_logic;
signal wdtick_cnt_16 : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal wdtick_cnt_17 : std_logic;
signal n20782 : std_logic;
signal wdtick_cnt_18 : std_logic;
signal n20783 : std_logic;
signal wdtick_cnt_19 : std_logic;
signal n20784 : std_logic;
signal wdtick_cnt_20 : std_logic;
signal n20785 : std_logic;
signal wdtick_cnt_21 : std_logic;
signal n20786 : std_logic;
signal wdtick_cnt_22 : std_logic;
signal n20787 : std_logic;
signal wdtick_cnt_23 : std_logic;
signal n20788 : std_logic;
signal n20789 : std_logic;
signal n49 : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal wdtick_cnt_24 : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal n12366 : std_logic;
signal n7_adj_1757 : std_logic;
signal \n2562_cascade_\ : std_logic;
signal n15378 : std_logic;
signal n8_adj_1782 : std_logic;
signal n12540 : std_logic;
signal n14_adj_1606 : std_logic;
signal n22238 : std_logic;
signal \n22240_cascade_\ : std_logic;
signal n23053 : std_logic;
signal \n11280_cascade_\ : std_logic;
signal \n12509_cascade_\ : std_logic;
signal comm_length_2 : std_logic;
signal comm_length_0 : std_logic;
signal buf_adcdata_vac_17 : std_logic;
signal n23486 : std_logic;
signal buf_adcdata_vdc_17 : std_logic;
signal \n46_cascade_\ : std_logic;
signal comm_test_buf_24_0 : std_logic;
signal comm_test_buf_24_8 : std_logic;
signal n14_adj_1662 : std_logic;
signal n4_adj_1749 : std_logic;
signal n12_adj_1684 : std_logic;
signal n14_adj_1608 : std_logic;
signal n13129 : std_logic;
signal \buf_cfgRTD_0\ : std_logic;
signal n22351 : std_logic;
signal \n4_adj_1709_cascade_\ : std_logic;
signal n35 : std_logic;
signal n12_adj_1802 : std_logic;
signal \comm_buf_1_7_N_559_3\ : std_logic;
signal comm_buf_1_3 : std_logic;
signal comm_buf_1_6 : std_logic;
signal comm_buf_1_0 : std_logic;
signal data_idxvec_14 : std_logic;
signal n22296 : std_logic;
signal data_idxvec_12 : std_logic;
signal n22499 : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal req_data_cnt_6 : std_logic;
signal \n23519_cascade_\ : std_logic;
signal n23291 : std_logic;
signal n111_adj_1726 : std_logic;
signal \n30_adj_1724_cascade_\ : std_logic;
signal \comm_buf_1_7_N_559_6\ : std_logic;
signal data_idxvec_6 : std_logic;
signal \n26_adj_1723_cascade_\ : std_logic;
signal n23516 : std_logic;
signal n23303 : std_logic;
signal n23555 : std_logic;
signal n18363 : std_logic;
signal buf_dds1_4 : std_logic;
signal \iac_raw_buf_N_823\ : std_logic;
signal data_cntvec_0 : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal n20622 : std_logic;
signal n20623 : std_logic;
signal data_cntvec_3 : std_logic;
signal n20624 : std_logic;
signal n20625 : std_logic;
signal n20626 : std_logic;
signal data_cntvec_6 : std_logic;
signal n20627 : std_logic;
signal n20628 : std_logic;
signal n20629 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal data_cntvec_8 : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal n20630 : std_logic;
signal data_cntvec_10 : std_logic;
signal n20631 : std_logic;
signal n20632 : std_logic;
signal data_cntvec_12 : std_logic;
signal n20633 : std_logic;
signal data_cntvec_13 : std_logic;
signal n20634 : std_logic;
signal n20635 : std_logic;
signal n20636 : std_logic;
signal data_cntvec_15 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal n12394 : std_logic;
signal n15431 : std_logic;
signal n23480 : std_logic;
signal \DDS_RNG_0\ : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal \n22183_cascade_\ : std_logic;
signal n22177 : std_logic;
signal n22180 : std_logic;
signal \n23462_cascade_\ : std_logic;
signal n23465 : std_logic;
signal data_idxvec_9 : std_logic;
signal data_cntvec_9 : std_logic;
signal buf_data_iac_17 : std_logic;
signal \n22184_cascade_\ : std_logic;
signal n22186 : std_logic;
signal n21997 : std_logic;
signal n14_adj_1656 : std_logic;
signal n13093 : std_logic;
signal buf_dds0_9 : std_logic;
signal dds_state_0 : std_logic;
signal dds_state_2 : std_logic;
signal dds_state_1 : std_logic;
signal \DDS_CS\ : std_logic;
signal \SIG_DDS.n9_adj_1490\ : std_logic;
signal buf_data_iac_23 : std_logic;
signal n22595 : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_840\ : std_logic;
signal \comm_spi.n24034\ : std_logic;
signal \comm_spi.n15352\ : std_logic;
signal \comm_spi.n15353\ : std_logic;
signal \comm_spi.n15357\ : std_logic;
signal \comm_spi.data_tx_7__N_874\ : std_logic;
signal \n22489_cascade_\ : std_logic;
signal \n20959_cascade_\ : std_logic;
signal n21883 : std_logic;
signal n19241 : std_logic;
signal n22033 : std_logic;
signal \n12064_cascade_\ : std_logic;
signal n21885 : std_logic;
signal \n22073_cascade_\ : std_logic;
signal flagcntwd : std_logic;
signal n12050 : std_logic;
signal n10_adj_1602 : std_logic;
signal comm_cmd_7 : std_logic;
signal n29 : std_logic;
signal n12951 : std_logic;
signal n9714 : std_logic;
signal n11_adj_1585 : std_logic;
signal n14_adj_1652 : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal n22487 : std_logic;
signal n21983 : std_logic;
signal n13171 : std_logic;
signal \n13171_cascade_\ : std_logic;
signal n22354 : std_logic;
signal n22353 : std_logic;
signal comm_length_1 : std_logic;
signal n4_adj_1745 : std_logic;
signal comm_index_1 : std_logic;
signal req_data_cnt_14 : std_logic;
signal data_cntvec_14 : std_logic;
signal n23 : std_logic;
signal n111 : std_logic;
signal n30_adj_1579 : std_logic;
signal \comm_buf_1_7_N_559_0\ : std_logic;
signal n21271 : std_logic;
signal n11258 : std_logic;
signal n22089 : std_logic;
signal n20318 : std_logic;
signal \n12_adj_1677_cascade_\ : std_logic;
signal \n12892_cascade_\ : std_logic;
signal \n37_cascade_\ : std_logic;
signal \n12761_cascade_\ : std_logic;
signal data_idxvec_5 : std_logic;
signal data_cntvec_5 : std_logic;
signal \n26_adj_1730_cascade_\ : std_logic;
signal req_data_cnt_5 : std_logic;
signal \n23336_cascade_\ : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal \n23339_cascade_\ : std_logic;
signal \n30_adj_1731_cascade_\ : std_logic;
signal n111_adj_1732 : std_logic;
signal \comm_buf_1_7_N_559_5_cascade_\ : std_logic;
signal n16_adj_1728 : std_logic;
signal buf_adcdata_iac_13 : std_logic;
signal n23354 : std_logic;
signal n23357 : std_logic;
signal data_idxvec_1 : std_logic;
signal data_cntvec_1 : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal req_data_cnt_1 : std_logic;
signal \n22142_cascade_\ : std_logic;
signal n22137 : std_logic;
signal \n23408_cascade_\ : std_logic;
signal \n23411_cascade_\ : std_logic;
signal n111_adj_1754 : std_logic;
signal \comm_buf_1_7_N_559_1_cascade_\ : std_logic;
signal comm_buf_1_1 : std_logic;
signal buf_data_iac_9 : std_logic;
signal n26_adj_1753 : std_logic;
signal n22143 : std_logic;
signal data_idxvec_4 : std_logic;
signal data_cntvec_4 : std_logic;
signal n22301 : std_logic;
signal \n26_adj_1735_cascade_\ : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal \n23318_cascade_\ : std_logic;
signal req_data_cnt_4 : std_logic;
signal n23441 : std_logic;
signal \n23321_cascade_\ : std_logic;
signal n111_adj_1737 : std_logic;
signal \n30_adj_1736_cascade_\ : std_logic;
signal \comm_buf_1_7_N_559_4_cascade_\ : std_logic;
signal data_idxvec_2 : std_logic;
signal data_cntvec_2 : std_logic;
signal buf_data_iac_10 : std_logic;
signal \n26_adj_1748_cascade_\ : std_logic;
signal \n22152_cascade_\ : std_logic;
signal n22149 : std_logic;
signal \n23444_cascade_\ : std_logic;
signal n22148 : std_logic;
signal n111_adj_1750 : std_logic;
signal \n23447_cascade_\ : std_logic;
signal \comm_buf_1_7_N_559_2_cascade_\ : std_logic;
signal comm_buf_1_2 : std_logic;
signal req_data_cnt_2 : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal n22151 : std_logic;
signal \SELIRNG1\ : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal buf_adcdata_iac_9 : std_logic;
signal n16_adj_1751 : std_logic;
signal n22136 : std_logic;
signal wdtick_flag : std_logic;
signal buf_control_0 : std_logic;
signal \CONT_SD\ : std_logic;
signal n8_adj_1605 : std_logic;
signal n7 : std_logic;
signal \data_index_9_N_236_0\ : std_logic;
signal buf_data_iac_20 : std_logic;
signal n22500 : std_logic;
signal \bfn_19_5_0_\ : std_logic;
signal \ADC_VDC.genclk.n20751\ : std_logic;
signal \ADC_VDC.genclk.n20752\ : std_logic;
signal \ADC_VDC.genclk.n20753\ : std_logic;
signal \ADC_VDC.genclk.n20754\ : std_logic;
signal \ADC_VDC.genclk.n20755\ : std_logic;
signal \ADC_VDC.genclk.n20756\ : std_logic;
signal \ADC_VDC.genclk.n20757\ : std_logic;
signal \ADC_VDC.genclk.n20758\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i0C_net\ : std_logic;
signal \bfn_19_6_0_\ : std_logic;
signal \ADC_VDC.genclk.n20759\ : std_logic;
signal \ADC_VDC.genclk.n20760\ : std_logic;
signal \ADC_VDC.genclk.n20761\ : std_logic;
signal \ADC_VDC.genclk.n20762\ : std_logic;
signal \ADC_VDC.genclk.n20763\ : std_logic;
signal \ADC_VDC.genclk.n20764\ : std_logic;
signal \ADC_VDC.genclk.n20765\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i8C_net\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal n20819 : std_logic;
signal n20820 : std_logic;
signal n20821 : std_logic;
signal n20822 : std_logic;
signal n20823 : std_logic;
signal n20824 : std_logic;
signal n20825 : std_logic;
signal \INVdds0_mclkcnt_i7_3792__i0C_net\ : std_logic;
signal n10 : std_logic;
signal dds0_mclkcnt_6 : std_logic;
signal \DDS_MCLK\ : std_logic;
signal \INVdds0_mclk_297C_net\ : std_logic;
signal \n6888_cascade_\ : std_logic;
signal n21865 : std_logic;
signal n21981 : std_logic;
signal n22027 : std_logic;
signal n22018 : std_logic;
signal dds0_mclkcnt_3 : std_logic;
signal dds0_mclkcnt_5 : std_logic;
signal dds0_mclkcnt_1 : std_logic;
signal dds0_mclkcnt_4 : std_logic;
signal dds0_mclkcnt_7 : std_logic;
signal dds0_mclkcnt_0 : std_logic;
signal \n12_adj_1685_cascade_\ : std_logic;
signal dds0_mclkcnt_2 : std_logic;
signal n21857 : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.n18536\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal n22330 : std_logic;
signal n22329 : std_logic;
signal n15261 : std_logic;
signal \n22321_cascade_\ : std_logic;
signal n14851 : std_logic;
signal n22352 : std_logic;
signal comm_index_2 : std_logic;
signal n21956 : std_logic;
signal n21862 : std_logic;
signal comm_index_0 : std_logic;
signal \n21862_cascade_\ : std_logic;
signal n30_adj_1720 : std_logic;
signal n21968 : std_logic;
signal \n22_adj_1725_cascade_\ : std_logic;
signal \n12677_cascade_\ : std_logic;
signal n21895 : std_logic;
signal buf_data_vac_8 : std_logic;
signal comm_rx_buf_0 : std_logic;
signal comm_buf_4_0 : std_logic;
signal buf_data_vac_15 : std_logic;
signal comm_buf_4_7 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal buf_data_vac_14 : std_logic;
signal comm_buf_4_6 : std_logic;
signal comm_rx_buf_5 : std_logic;
signal buf_data_vac_13 : std_logic;
signal comm_buf_4_5 : std_logic;
signal comm_rx_buf_4 : std_logic;
signal buf_data_vac_12 : std_logic;
signal comm_buf_4_4 : std_logic;
signal buf_data_vac_11 : std_logic;
signal comm_buf_4_3 : std_logic;
signal comm_rx_buf_2 : std_logic;
signal buf_data_vac_10 : std_logic;
signal comm_buf_4_2 : std_logic;
signal comm_rx_buf_1 : std_logic;
signal buf_data_vac_9 : std_logic;
signal comm_buf_4_1 : std_logic;
signal n12892 : std_logic;
signal n15510 : std_logic;
signal data_idxvec_7 : std_logic;
signal data_cntvec_7 : std_logic;
signal buf_data_iac_15 : std_logic;
signal \n26_adj_1716_cascade_\ : std_logic;
signal \n22263_cascade_\ : std_logic;
signal n22272 : std_logic;
signal \n23420_cascade_\ : std_logic;
signal n22271 : std_logic;
signal n111_adj_1719 : std_logic;
signal \n23423_cascade_\ : std_logic;
signal comm_rx_buf_7 : std_logic;
signal \comm_buf_1_7_N_559_7_cascade_\ : std_logic;
signal comm_buf_1_7 : std_logic;
signal n12761 : std_logic;
signal n15489 : std_logic;
signal n18955 : std_logic;
signal n22356 : std_logic;
signal buf_dds0_13 : std_logic;
signal n23348 : std_logic;
signal req_data_cnt_7 : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal n22262 : std_logic;
signal buf_data_iac_14 : std_logic;
signal n22391 : std_logic;
signal n12509 : std_logic;
signal n14_adj_1660 : std_logic;
signal buf_dds1_13 : std_logic;
signal comm_buf_1_5 : std_logic;
signal data_index_5 : std_logic;
signal n9324 : std_logic;
signal n8_adj_1623 : std_logic;
signal \n8_adj_1623_cascade_\ : std_logic;
signal n7_adj_1622 : std_logic;
signal \data_index_9_N_236_5\ : std_logic;
signal n21966 : std_logic;
signal trig_dds1 : std_logic;
signal n21920 : std_logic;
signal \n22399_cascade_\ : std_logic;
signal n40_adj_1689 : std_logic;
signal data_idxvec_11 : std_logic;
signal data_cntvec_11 : std_logic;
signal comm_buf_1_4 : std_logic;
signal n14_adj_1611 : std_logic;
signal n14_adj_1654 : std_logic;
signal \INVADC_VDC.genclk.div_state_i1C_net\ : std_logic;
signal \ADC_VDC.genclk.n6\ : std_logic;
signal \ADC_VDC.genclk.t0on_6\ : std_logic;
signal \ADC_VDC.genclk.t0on_1\ : std_logic;
signal \ADC_VDC.genclk.t0on_4\ : std_logic;
signal \ADC_VDC.genclk.t0on_0\ : std_logic;
signal \ADC_VDC.genclk.n22308_cascade_\ : std_logic;
signal \ADC_VDC.genclk.t0on_12\ : std_logic;
signal \ADC_VDC.genclk.t0on_2\ : std_logic;
signal \ADC_VDC.genclk.t0on_7\ : std_logic;
signal \ADC_VDC.genclk.t0on_10\ : std_logic;
signal \ADC_VDC.genclk.n27_adj_1483\ : std_logic;
signal \ADC_VDC.genclk.t0on_14\ : std_logic;
signal \ADC_VDC.genclk.t0on_9\ : std_logic;
signal \ADC_VDC.genclk.t0on_15\ : std_logic;
signal \ADC_VDC.genclk.t0on_11\ : std_logic;
signal \ADC_VDC.genclk.n28_adj_1481\ : std_logic;
signal \ADC_VDC.genclk.t0on_13\ : std_logic;
signal \ADC_VDC.genclk.t0on_3\ : std_logic;
signal \ADC_VDC.genclk.t0on_5\ : std_logic;
signal \ADC_VDC.genclk.t0on_8\ : std_logic;
signal \ADC_VDC.genclk.n26_adj_1482\ : std_logic;
signal \ADC_VDC.genclk.div_state_1__N_1480\ : std_logic;
signal comm_clear : std_logic;
signal buf_data_iac_18 : std_logic;
signal n22170 : std_logic;
signal n12035 : std_logic;
signal n7_adj_1687 : std_logic;
signal \comm_state_3_N_484_3\ : std_logic;
signal n1373 : std_logic;
signal \n2_cascade_\ : std_logic;
signal n23342 : std_logic;
signal n9837 : std_logic;
signal \n23345_cascade_\ : std_logic;
signal n8_adj_1659 : std_logic;
signal n2562 : std_logic;
signal n22339 : std_logic;
signal \n22340_cascade_\ : std_logic;
signal n14_adj_1593 : std_logic;
signal n5 : std_logic;
signal \n9725_cascade_\ : std_logic;
signal n4 : std_logic;
signal n22492 : std_logic;
signal \n6_adj_1657_cascade_\ : std_logic;
signal \n26_adj_1597_cascade_\ : std_logic;
signal n18_adj_1595 : std_logic;
signal n21908 : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal comm_data_vld : std_logic;
signal n4_adj_1718 : std_logic;
signal req_data_cnt_11 : std_logic;
signal n112_adj_1777 : std_logic;
signal \comm_buf_0_7_N_543_5\ : std_logic;
signal comm_cmd_5 : std_logic;
signal comm_cmd_4 : std_logic;
signal n22365 : std_logic;
signal \n22364_cascade_\ : std_logic;
signal n48 : std_logic;
signal \n22370_cascade_\ : std_logic;
signal n7148 : std_logic;
signal n22368 : std_logic;
signal n9_adj_1507 : std_logic;
signal n23387 : std_logic;
signal n23351 : std_logic;
signal n23495 : std_logic;
signal buf_data_iac_19 : std_logic;
signal n22642 : std_logic;
signal n23_adj_1791 : std_logic;
signal n23501 : std_logic;
signal \n23459_cascade_\ : std_logic;
signal n112_adj_1795 : std_logic;
signal \n30_adj_1793_cascade_\ : std_logic;
signal comm_cmd_6 : std_logic;
signal data_idxvec_13 : std_logic;
signal buf_data_iac_21 : std_logic;
signal \n28_adj_1775_cascade_\ : std_logic;
signal comm_cmd_3 : std_logic;
signal n23492 : std_logic;
signal n23_adj_1773 : std_logic;
signal req_data_cnt_13 : std_logic;
signal n25_adj_1774 : std_logic;
signal comm_cmd_1 : std_logic;
signal comm_cmd_2 : std_logic;
signal n22316 : std_logic;
signal n26_adj_1792 : std_logic;
signal n23456 : std_logic;
signal buf_data_iac_13 : std_logic;
signal n22313 : std_logic;
signal buf_data_iac_11 : std_logic;
signal n22300 : std_logic;
signal buf_data_iac_8 : std_logic;
signal comm_cmd_0 : std_logic;
signal n22649 : std_logic;
signal \ADC_VDC.genclk.n26\ : std_logic;
signal \ADC_VDC.genclk.n22305_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n27\ : std_logic;
signal \ADC_VDC.genclk.n22303\ : std_logic;
signal \ADC_VDC.genclk.div_state_1\ : std_logic;
signal \ADC_VDC.genclk.n22303_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n22302\ : std_logic;
signal \ADC_VDC.genclk.div_state_0\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.n28\ : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal comm_state_2 : std_logic;
signal comm_state_3 : std_logic;
signal n12966 : std_logic;
signal comm_state_0 : std_logic;
signal n12045 : std_logic;
signal comm_rx_buf_3 : std_logic;
signal comm_state_1 : std_logic;
signal \comm_buf_0_7_N_543_3\ : std_logic;
signal comm_buf_0_3 : std_logic;
signal \clk_32MHz\ : std_logic;
signal n12677 : std_logic;
signal n15482 : std_logic;
signal \ADC_VDC.genclk.t0off_0\ : std_logic;
signal \bfn_23_5_0_\ : std_logic;
signal \ADC_VDC.genclk.t0off_1\ : std_logic;
signal \ADC_VDC.genclk.n20736\ : std_logic;
signal \ADC_VDC.genclk.t0off_2\ : std_logic;
signal \ADC_VDC.genclk.n20737\ : std_logic;
signal \ADC_VDC.genclk.t0off_3\ : std_logic;
signal \ADC_VDC.genclk.n20738\ : std_logic;
signal \ADC_VDC.genclk.t0off_4\ : std_logic;
signal \ADC_VDC.genclk.n20739\ : std_logic;
signal \ADC_VDC.genclk.t0off_5\ : std_logic;
signal \ADC_VDC.genclk.n20740\ : std_logic;
signal \ADC_VDC.genclk.t0off_6\ : std_logic;
signal \ADC_VDC.genclk.n20741\ : std_logic;
signal \ADC_VDC.genclk.t0off_7\ : std_logic;
signal \ADC_VDC.genclk.n20742\ : std_logic;
signal \ADC_VDC.genclk.n20743\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.t0off_8\ : std_logic;
signal \bfn_23_6_0_\ : std_logic;
signal \ADC_VDC.genclk.t0off_9\ : std_logic;
signal \ADC_VDC.genclk.n20744\ : std_logic;
signal \ADC_VDC.genclk.t0off_10\ : std_logic;
signal \ADC_VDC.genclk.n20745\ : std_logic;
signal \ADC_VDC.genclk.t0off_11\ : std_logic;
signal \ADC_VDC.genclk.n20746\ : std_logic;
signal \ADC_VDC.genclk.t0off_12\ : std_logic;
signal \ADC_VDC.genclk.n20747\ : std_logic;
signal \ADC_VDC.genclk.t0off_13\ : std_logic;
signal \ADC_VDC.genclk.n20748\ : std_logic;
signal \ADC_VDC.genclk.t0off_14\ : std_logic;
signal \ADC_VDC.genclk.n20749\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ADC_VDC.genclk.n20750\ : std_logic;
signal \ADC_VDC.genclk.t0off_15\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.n12361\ : std_logic;
signal \ADC_VDC.genclk.n15418\ : std_logic;

signal \VAC_DRDY_wire\ : std_logic;
signal \IAC_FLT1_wire\ : std_logic;
signal \DDS_SCK_wire\ : std_logic;
signal \ICE_IOR_166_wire\ : std_logic;
signal \ICE_IOR_119_wire\ : std_logic;
signal \DDS_MOSI_wire\ : std_logic;
signal \VAC_MISO_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \ICE_IOR_146_wire\ : std_logic;
signal \VDC_CLK_wire\ : std_logic;
signal \ICE_IOT_222_wire\ : std_logic;
signal \IAC_CS_wire\ : std_logic;
signal \ICE_IOL_18B_wire\ : std_logic;
signal \ICE_IOL_13A_wire\ : std_logic;
signal \ICE_IOB_81_wire\ : std_logic;
signal \VAC_OSR1_wire\ : std_logic;
signal \IAC_MOSI_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \ICE_IOL_4B_wire\ : std_logic;
signal \ICE_IOB_94_wire\ : std_logic;
signal \VAC_CS_wire\ : std_logic;
signal \VAC_CLK_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \ICE_IOR_167_wire\ : std_logic;
signal \ICE_IOR_118_wire\ : std_logic;
signal \RTD_SDO_wire\ : std_logic;
signal \IAC_OSR0_wire\ : std_logic;
signal \VDC_SCLK_wire\ : std_logic;
signal \VAC_FLT1_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_IOR_165_wire\ : std_logic;
signal \ICE_IOR_147_wire\ : std_logic;
signal \ICE_IOL_14A_wire\ : std_logic;
signal \ICE_IOL_13B_wire\ : std_logic;
signal \ICE_IOB_91_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_RNG_0_wire\ : std_logic;
signal \VDC_RNG0_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \ICE_IOR_152_wire\ : std_logic;
signal \ICE_IOL_12A_wire\ : std_logic;
signal \RTD_DRDY_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_IOT_177_wire\ : std_logic;
signal \ICE_IOR_141_wire\ : std_logic;
signal \ICE_IOB_80_wire\ : std_logic;
signal \ICE_IOB_102_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \IAC_MISO_wire\ : std_logic;
signal \VAC_OSR0_wire\ : std_logic;
signal \VAC_MOSI_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \ICE_IOR_148_wire\ : std_logic;
signal \STAT_COMM_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \ICE_IOR_161_wire\ : std_logic;
signal \ICE_IOB_95_wire\ : std_logic;
signal \ICE_IOB_82_wire\ : std_logic;
signal \ICE_IOB_104_wire\ : std_logic;
signal \IAC_CLK_wire\ : std_logic;
signal \DDS_CS_wire\ : std_logic;
signal \SELIRNG0_wire\ : std_logic;
signal \RTD_SDI_wire\ : std_logic;
signal \ICE_IOT_221_wire\ : std_logic;
signal \ICE_IOT_197_wire\ : std_logic;
signal \DDS_MCLK_wire\ : std_logic;
signal \RTD_SCLK_wire\ : std_logic;
signal \RTD_CS_wire\ : std_logic;
signal \ICE_IOR_137_wire\ : std_logic;
signal \IAC_OSR1_wire\ : std_logic;
signal \VAC_FLT0_wire\ : std_logic;
signal \ICE_IOR_144_wire\ : std_logic;
signal \ICE_IOR_128_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \IAC_SCLK_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \ICE_IOR_139_wire\ : std_logic;
signal \ICE_IOL_4A_wire\ : std_logic;
signal \VAC_SCLK_wire\ : std_logic;
signal \THERMOSTAT_wire\ : std_logic;
signal \ICE_IOR_164_wire\ : std_logic;
signal \ICE_IOB_103_wire\ : std_logic;
signal \AMPV_POW_wire\ : std_logic;
signal \VDC_SDO_wire\ : std_logic;
signal \ICE_IOT_174_wire\ : std_logic;
signal \ICE_IOR_140_wire\ : std_logic;
signal \ICE_IOB_96_wire\ : std_logic;
signal \CONT_SD_wire\ : std_logic;
signal \AC_ADC_SYNC_wire\ : std_logic;
signal \SELIRNG1_wire\ : std_logic;
signal \ICE_IOL_12B_wire\ : std_logic;
signal \ICE_IOR_160_wire\ : std_logic;
signal \ICE_IOR_136_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_IOT_198_wire\ : std_logic;
signal \ICE_IOT_173_wire\ : std_logic;
signal \IAC_DRDY_wire\ : std_logic;
signal \ICE_IOT_178_wire\ : std_logic;
signal \ICE_IOR_138_wire\ : std_logic;
signal \ICE_IOR_120_wire\ : std_logic;
signal \IAC_FLT0_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \VAC_DRDY_wire\ <= VAC_DRDY;
    IAC_FLT1 <= \IAC_FLT1_wire\;
    DDS_SCK <= \DDS_SCK_wire\;
    \ICE_IOR_166_wire\ <= ICE_IOR_166;
    \ICE_IOR_119_wire\ <= ICE_IOR_119;
    DDS_MOSI <= \DDS_MOSI_wire\;
    \VAC_MISO_wire\ <= VAC_MISO;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    \ICE_IOR_146_wire\ <= ICE_IOR_146;
    VDC_CLK <= \VDC_CLK_wire\;
    \ICE_IOT_222_wire\ <= ICE_IOT_222;
    IAC_CS <= \IAC_CS_wire\;
    \ICE_IOL_18B_wire\ <= ICE_IOL_18B;
    \ICE_IOL_13A_wire\ <= ICE_IOL_13A;
    \ICE_IOB_81_wire\ <= ICE_IOB_81;
    VAC_OSR1 <= \VAC_OSR1_wire\;
    IAC_MOSI <= \IAC_MOSI_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    \ICE_IOL_4B_wire\ <= ICE_IOL_4B;
    \ICE_IOB_94_wire\ <= ICE_IOB_94;
    VAC_CS <= \VAC_CS_wire\;
    VAC_CLK <= \VAC_CLK_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    \ICE_IOR_167_wire\ <= ICE_IOR_167;
    \ICE_IOR_118_wire\ <= ICE_IOR_118;
    \RTD_SDO_wire\ <= RTD_SDO;
    IAC_OSR0 <= \IAC_OSR0_wire\;
    VDC_SCLK <= \VDC_SCLK_wire\;
    VAC_FLT1 <= \VAC_FLT1_wire\;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_IOR_165_wire\ <= ICE_IOR_165;
    \ICE_IOR_147_wire\ <= ICE_IOR_147;
    \ICE_IOL_14A_wire\ <= ICE_IOL_14A;
    \ICE_IOL_13B_wire\ <= ICE_IOL_13B;
    \ICE_IOB_91_wire\ <= ICE_IOB_91;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_RNG_0 <= \DDS_RNG_0_wire\;
    VDC_RNG0 <= \VDC_RNG0_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    \ICE_IOR_152_wire\ <= ICE_IOR_152;
    \ICE_IOL_12A_wire\ <= ICE_IOL_12A;
    \RTD_DRDY_wire\ <= RTD_DRDY;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_IOT_177_wire\ <= ICE_IOT_177;
    \ICE_IOR_141_wire\ <= ICE_IOR_141;
    \ICE_IOB_80_wire\ <= ICE_IOB_80;
    \ICE_IOB_102_wire\ <= ICE_IOB_102;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    \IAC_MISO_wire\ <= IAC_MISO;
    VAC_OSR0 <= \VAC_OSR0_wire\;
    VAC_MOSI <= \VAC_MOSI_wire\;
    TEST_LED <= \TEST_LED_wire\;
    \ICE_IOR_148_wire\ <= ICE_IOR_148;
    STAT_COMM <= \STAT_COMM_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    \ICE_IOR_161_wire\ <= ICE_IOR_161;
    \ICE_IOB_95_wire\ <= ICE_IOB_95;
    \ICE_IOB_82_wire\ <= ICE_IOB_82;
    \ICE_IOB_104_wire\ <= ICE_IOB_104;
    IAC_CLK <= \IAC_CLK_wire\;
    DDS_CS <= \DDS_CS_wire\;
    SELIRNG0 <= \SELIRNG0_wire\;
    RTD_SDI <= \RTD_SDI_wire\;
    \ICE_IOT_221_wire\ <= ICE_IOT_221;
    \ICE_IOT_197_wire\ <= ICE_IOT_197;
    DDS_MCLK <= \DDS_MCLK_wire\;
    RTD_SCLK <= \RTD_SCLK_wire\;
    RTD_CS <= \RTD_CS_wire\;
    \ICE_IOR_137_wire\ <= ICE_IOR_137;
    IAC_OSR1 <= \IAC_OSR1_wire\;
    VAC_FLT0 <= \VAC_FLT0_wire\;
    \ICE_IOR_144_wire\ <= ICE_IOR_144;
    \ICE_IOR_128_wire\ <= ICE_IOR_128;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    IAC_SCLK <= \IAC_SCLK_wire\;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    \ICE_IOR_139_wire\ <= ICE_IOR_139;
    \ICE_IOL_4A_wire\ <= ICE_IOL_4A;
    VAC_SCLK <= \VAC_SCLK_wire\;
    \THERMOSTAT_wire\ <= THERMOSTAT;
    \ICE_IOR_164_wire\ <= ICE_IOR_164;
    \ICE_IOB_103_wire\ <= ICE_IOB_103;
    AMPV_POW <= \AMPV_POW_wire\;
    \VDC_SDO_wire\ <= VDC_SDO;
    \ICE_IOT_174_wire\ <= ICE_IOT_174;
    \ICE_IOR_140_wire\ <= ICE_IOR_140;
    \ICE_IOB_96_wire\ <= ICE_IOB_96;
    CONT_SD <= \CONT_SD_wire\;
    AC_ADC_SYNC <= \AC_ADC_SYNC_wire\;
    SELIRNG1 <= \SELIRNG1_wire\;
    \ICE_IOL_12B_wire\ <= ICE_IOL_12B;
    \ICE_IOR_160_wire\ <= ICE_IOR_160;
    \ICE_IOR_136_wire\ <= ICE_IOR_136;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_IOT_198_wire\ <= ICE_IOT_198;
    \ICE_IOT_173_wire\ <= ICE_IOT_173;
    \IAC_DRDY_wire\ <= IAC_DRDY;
    \ICE_IOT_178_wire\ <= ICE_IOT_178;
    \ICE_IOR_138_wire\ <= ICE_IOR_138;
    \ICE_IOR_120_wire\ <= ICE_IOR_120;
    IAC_FLT0 <= \IAC_FLT0_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data_iac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(13);
    buf_data_vac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(9);
    buf_data_iac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(5);
    buf_data_vac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ <= '0'&\N__44452\&\N__42274\&\N__44878\&\N__45073\&\N__56338\&\N__43771\&\N__39061\&\N__41731\&\N__40135\&\N__53098\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ <= '0'&\N__29899\&\N__30007\&\N__30115\&\N__30214\&\N__29152\&\N__29260\&\N__29365\&\N__29473\&\N__29584\&\N__29686\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ <= '0'&'0'&\N__28003\&'0'&'0'&'0'&\N__27841\&'0'&'0'&'0'&\N__30610\&'0'&'0'&'0'&\N__31495\&'0';
    buf_data_iac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(13);
    buf_data_vac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(9);
    buf_data_iac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(5);
    buf_data_vac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ <= '0'&\N__44412\&\N__42231\&\N__44835\&\N__45030\&\N__56289\&\N__43725\&\N__39018\&\N__41685\&\N__40092\&\N__53055\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ <= '0'&\N__29865\&\N__29970\&\N__30078\&\N__30180\&\N__29115\&\N__29223\&\N__29328\&\N__29439\&\N__29553\&\N__29649\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ <= '0'&'0'&\N__52720\&'0'&'0'&'0'&\N__23878\&'0'&'0'&'0'&\N__46956\&'0'&'0'&'0'&\N__25300\&'0';
    buf_data_iac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(13);
    buf_data_vac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(9);
    buf_data_iac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(5);
    buf_data_vac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ <= '0'&\N__44470\&\N__42292\&\N__44896\&\N__45091\&\N__56356\&\N__43789\&\N__39079\&\N__41749\&\N__40153\&\N__53116\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ <= '0'&\N__29917\&\N__30025\&\N__30133\&\N__30232\&\N__29170\&\N__29278\&\N__29383\&\N__29491\&\N__29602\&\N__29704\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ <= '0'&'0'&\N__38623\&'0'&'0'&'0'&\N__31210\&'0'&'0'&'0'&\N__37171\&'0'&'0'&'0'&\N__25459\&'0';
    buf_data_iac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(13);
    buf_data_vac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(9);
    buf_data_iac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(5);
    buf_data_vac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ <= '0'&\N__44424\&\N__42243\&\N__44847\&\N__45042\&\N__56301\&\N__43737\&\N__39030\&\N__41697\&\N__40104\&\N__53067\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ <= '0'&\N__29875\&\N__29982\&\N__30090\&\N__30190\&\N__29127\&\N__29235\&\N__29340\&\N__29449\&\N__29560\&\N__29661\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ <= '0'&'0'&\N__44229\&'0'&'0'&'0'&\N__41230\&'0'&'0'&'0'&\N__42076\&'0'&'0'&'0'&\N__25087\&'0';
    buf_data_iac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(13);
    buf_data_vac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(9);
    buf_data_iac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(5);
    buf_data_vac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ <= '0'&\N__44476\&\N__42298\&\N__44902\&\N__45097\&\N__56362\&\N__43795\&\N__39085\&\N__41755\&\N__40159\&\N__53122\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ <= '0'&\N__29923\&\N__30031\&\N__30139\&\N__30238\&\N__29176\&\N__29284\&\N__29389\&\N__29497\&\N__29608\&\N__29710\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ <= '0'&'0'&\N__25402\&'0'&'0'&'0'&\N__23254\&'0'&'0'&'0'&\N__31690\&'0'&'0'&'0'&\N__23104\&'0';
    buf_data_iac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(13);
    buf_data_vac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(9);
    buf_data_iac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(5);
    buf_data_vac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ <= '0'&\N__44434\&\N__42255\&\N__44859\&\N__45054\&\N__56313\&\N__43749\&\N__39042\&\N__41709\&\N__40116\&\N__53079\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ <= '0'&\N__29881\&\N__29989\&\N__30097\&\N__30196\&\N__29134\&\N__29242\&\N__29347\&\N__29455\&\N__29566\&\N__29668\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ <= '0'&'0'&\N__52341\&'0'&'0'&'0'&\N__38050\&'0'&'0'&'0'&\N__36985\&'0'&'0'&'0'&\N__30928\&'0';
    buf_data_iac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(13);
    buf_data_vac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(9);
    buf_data_iac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(5);
    buf_data_vac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ <= '0'&\N__44421\&\N__42246\&\N__44850\&\N__45045\&\N__56316\&\N__43746\&\N__39033\&\N__41706\&\N__40107\&\N__53070\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ <= '0'&\N__29862\&\N__29973\&\N__30081\&\N__30177\&\N__29118\&\N__29226\&\N__29331\&\N__29436\&\N__29544\&\N__29652\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ <= '0'&'0'&\N__22165\&'0'&'0'&'0'&\N__22930\&'0'&'0'&'0'&\N__21961\&'0'&'0'&'0'&\N__21562\&'0';
    buf_data_iac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(13);
    buf_data_vac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(9);
    buf_data_iac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(5);
    buf_data_vac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ <= '0'&\N__44440\&\N__42262\&\N__44866\&\N__45061\&\N__56325\&\N__43759\&\N__39049\&\N__41719\&\N__40123\&\N__53086\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ <= '0'&\N__29887\&\N__29995\&\N__30103\&\N__30202\&\N__29140\&\N__29248\&\N__29353\&\N__29461\&\N__29572\&\N__29674\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ <= '0'&'0'&\N__46924\&'0'&'0'&'0'&\N__24232\&'0'&'0'&'0'&\N__41310\&'0'&'0'&'0'&\N__28675\&'0';
    buf_data_iac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(13);
    buf_data_vac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(9);
    buf_data_iac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(5);
    buf_data_vac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ <= '0'&\N__44433\&\N__42258\&\N__44862\&\N__45057\&\N__56328\&\N__43758\&\N__39045\&\N__41718\&\N__40119\&\N__53082\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ <= '0'&\N__29874\&\N__29985\&\N__30093\&\N__30189\&\N__29130\&\N__29238\&\N__29343\&\N__29448\&\N__29556\&\N__29664\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ <= '0'&'0'&\N__22048\&'0'&'0'&'0'&\N__21988\&'0'&'0'&'0'&\N__22069\&'0'&'0'&'0'&\N__21865\&'0';
    buf_data_iac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(13);
    buf_data_vac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(9);
    buf_data_iac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(5);
    buf_data_vac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ <= '0'&\N__44464\&\N__42286\&\N__44890\&\N__45085\&\N__56350\&\N__43783\&\N__39073\&\N__41743\&\N__40147\&\N__53110\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ <= '0'&\N__29911\&\N__30019\&\N__30127\&\N__30226\&\N__29164\&\N__29272\&\N__29377\&\N__29485\&\N__29596\&\N__29698\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ <= '0'&'0'&\N__33700\&'0'&'0'&'0'&\N__33655\&'0'&'0'&'0'&\N__36067\&'0'&'0'&'0'&\N__35458\&'0';
    buf_data_iac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(13);
    buf_data_vac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(9);
    buf_data_iac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(5);
    buf_data_vac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ <= '0'&\N__44446\&\N__42268\&\N__44872\&\N__45067\&\N__56332\&\N__43765\&\N__39055\&\N__41725\&\N__40129\&\N__53092\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ <= '0'&\N__29893\&\N__30001\&\N__30109\&\N__30208\&\N__29146\&\N__29254\&\N__29359\&\N__29467\&\N__29578\&\N__29680\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ <= '0'&'0'&\N__30271\&'0'&'0'&'0'&\N__48613\&'0'&'0'&'0'&\N__34390\&'0'&'0'&'0'&\N__43516\&'0';
    buf_data_iac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(13);
    buf_data_vac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(9);
    buf_data_iac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(5);
    buf_data_vac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ <= '0'&\N__44458\&\N__42280\&\N__44884\&\N__45079\&\N__56344\&\N__43777\&\N__39067\&\N__41737\&\N__40141\&\N__53104\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ <= '0'&\N__29905\&\N__30013\&\N__30121\&\N__30220\&\N__29158\&\N__29266\&\N__29371\&\N__29479\&\N__29590\&\N__29692\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ <= '0'&'0'&\N__36094\&'0'&'0'&'0'&\N__33610\&'0'&'0'&'0'&\N__38098\&'0'&'0'&'0'&\N__37882\&'0';

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__21256\,
            RESETB => \N__64855\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \DDS_MCLK1\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \iac_raw_buf_vac_raw_buf_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61922\,
            RE => \N__64829\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            WE => \N__34523\
        );

    \iac_raw_buf_vac_raw_buf_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__62013\,
            RE => \N__64873\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            WE => \N__34522\
        );

    \iac_raw_buf_vac_raw_buf_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61852\,
            RE => \N__64824\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            WE => \N__34536\
        );

    \iac_raw_buf_vac_raw_buf_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__62010\,
            RE => \N__64869\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            WE => \N__34499\
        );

    \iac_raw_buf_vac_raw_buf_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61837\,
            RE => \N__64856\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            WE => \N__34540\
        );

    \iac_raw_buf_vac_raw_buf_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__62003\,
            RE => \N__64868\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            WE => \N__34498\
        );

    \iac_raw_buf_vac_raw_buf_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61881\,
            RE => \N__64617\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            WE => \N__34518\
        );

    \iac_raw_buf_vac_raw_buf_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61988\,
            RE => \N__64858\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            WE => \N__34503\
        );

    \iac_raw_buf_vac_raw_buf_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61859\,
            RE => \N__64616\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            WE => \N__34534\
        );

    \iac_raw_buf_vac_raw_buf_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61867\,
            RE => \N__64823\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            WE => \N__34535\
        );

    \iac_raw_buf_vac_raw_buf_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61959\,
            RE => \N__64857\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            WE => \N__34504\
        );

    \iac_raw_buf_vac_raw_buf_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__61892\,
            RE => \N__64828\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            WE => \N__34524\
        );

    \ipInertedIOPad_VAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65921\,
            DIN => \N__65920\,
            DOUT => \N__65919\,
            PACKAGEPIN => \VAC_DRDY_wire\
        );

    \ipInertedIOPad_VAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65921\,
            PADOUT => \N__65920\,
            PADIN => \N__65919\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65912\,
            DIN => \N__65911\,
            DOUT => \N__65910\,
            PACKAGEPIN => \IAC_FLT1_wire\
        );

    \ipInertedIOPad_IAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65912\,
            PADOUT => \N__65911\,
            PADIN => \N__65910\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29809\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65903\,
            DIN => \N__65902\,
            DOUT => \N__65901\,
            PACKAGEPIN => \DDS_SCK_wire\
        );

    \ipInertedIOPad_DDS_SCK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65903\,
            PADOUT => \N__65902\,
            PADIN => \N__65901\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__47614\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_166_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65894\,
            DIN => \N__65893\,
            DOUT => \N__65892\,
            PACKAGEPIN => \ICE_IOR_166_wire\
        );

    \ipInertedIOPad_ICE_IOR_166_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65894\,
            PADOUT => \N__65893\,
            PADIN => \N__65892\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_119_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65885\,
            DIN => \N__65884\,
            DOUT => \N__65883\,
            PACKAGEPIN => \ICE_IOR_119_wire\
        );

    \ipInertedIOPad_ICE_IOR_119_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65885\,
            PADOUT => \N__65884\,
            PADIN => \N__65883\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65876\,
            DIN => \N__65875\,
            DOUT => \N__65874\,
            PACKAGEPIN => \DDS_MOSI_wire\
        );

    \ipInertedIOPad_DDS_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65876\,
            PADOUT => \N__65875\,
            PADIN => \N__65874\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__40024\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65867\,
            DIN => \N__65866\,
            DOUT => \N__65865\,
            PACKAGEPIN => \VAC_MISO_wire\
        );

    \ipInertedIOPad_VAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65867\,
            PADOUT => \N__65866\,
            PADIN => \N__65865\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65858\,
            DIN => \N__65857\,
            DOUT => \N__65856\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65858\,
            PADOUT => \N__65857\,
            PADIN => \N__65856\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24289\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_146_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65849\,
            DIN => \N__65848\,
            DOUT => \N__65847\,
            PACKAGEPIN => \ICE_IOR_146_wire\
        );

    \ipInertedIOPad_ICE_IOR_146_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65849\,
            PADOUT => \N__65848\,
            PADIN => \N__65847\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65840\,
            DIN => \N__65839\,
            DOUT => \N__65838\,
            PACKAGEPIN => \VDC_CLK_wire\
        );

    \ipInertedIOPad_VDC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65840\,
            PADOUT => \N__65839\,
            PADIN => \N__65838\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42760\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_222_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65831\,
            DIN => \N__65830\,
            DOUT => \N__65829\,
            PACKAGEPIN => \ICE_IOT_222_wire\
        );

    \ipInertedIOPad_ICE_IOT_222_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65831\,
            PADOUT => \N__65830\,
            PADIN => \N__65829\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65822\,
            DIN => \N__65821\,
            DOUT => \N__65820\,
            PACKAGEPIN => \IAC_CS_wire\
        );

    \ipInertedIOPad_IAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65822\,
            PADOUT => \N__65821\,
            PADIN => \N__65820\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25771\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_18B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65813\,
            DIN => \N__65812\,
            DOUT => \N__65811\,
            PACKAGEPIN => \ICE_IOL_18B_wire\
        );

    \ipInertedIOPad_ICE_IOL_18B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65813\,
            PADOUT => \N__65812\,
            PADIN => \N__65811\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65804\,
            DIN => \N__65803\,
            DOUT => \N__65802\,
            PACKAGEPIN => \ICE_IOL_13A_wire\
        );

    \ipInertedIOPad_ICE_IOL_13A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65804\,
            PADOUT => \N__65803\,
            PADIN => \N__65802\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_81_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65795\,
            DIN => \N__65794\,
            DOUT => \N__65793\,
            PACKAGEPIN => \ICE_IOB_81_wire\
        );

    \ipInertedIOPad_ICE_IOB_81_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65795\,
            PADOUT => \N__65794\,
            PADIN => \N__65793\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65786\,
            DIN => \N__65785\,
            DOUT => \N__65784\,
            PACKAGEPIN => \VAC_OSR1_wire\
        );

    \ipInertedIOPad_VAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65786\,
            PADOUT => \N__65785\,
            PADIN => \N__65784\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__38668\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65777\,
            DIN => \N__65776\,
            DOUT => \N__65775\,
            PACKAGEPIN => \IAC_MOSI_wire\
        );

    \ipInertedIOPad_IAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65777\,
            PADOUT => \N__65776\,
            PADIN => \N__65775\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65768\,
            DIN => \N__65767\,
            DOUT => \N__65766\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65768\,
            PADOUT => \N__65767\,
            PADIN => \N__65766\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21658\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65759\,
            DIN => \N__65758\,
            DOUT => \N__65757\,
            PACKAGEPIN => \ICE_IOL_4B_wire\
        );

    \ipInertedIOPad_ICE_IOL_4B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65759\,
            PADOUT => \N__65758\,
            PADIN => \N__65757\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_94_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65750\,
            DIN => \N__65749\,
            DOUT => \N__65748\,
            PACKAGEPIN => \ICE_IOB_94_wire\
        );

    \ipInertedIOPad_ICE_IOB_94_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65750\,
            PADOUT => \N__65749\,
            PADIN => \N__65748\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65741\,
            DIN => \N__65740\,
            DOUT => \N__65739\,
            PACKAGEPIN => \VAC_CS_wire\
        );

    \ipInertedIOPad_VAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65741\,
            PADOUT => \N__65740\,
            PADIN => \N__65739\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21352\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65732\,
            DIN => \N__65731\,
            DOUT => \N__65730\,
            PACKAGEPIN => \VAC_CLK_wire\
        );

    \ipInertedIOPad_VAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65732\,
            PADOUT => \N__65731\,
            PADIN => \N__65730\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26026\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65723\,
            DIN => \N__65722\,
            DOUT => \N__65721\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65723\,
            PADOUT => \N__65722\,
            PADIN => \N__65721\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_167_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65714\,
            DIN => \N__65713\,
            DOUT => \N__65712\,
            PACKAGEPIN => \ICE_IOR_167_wire\
        );

    \ipInertedIOPad_ICE_IOR_167_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65714\,
            PADOUT => \N__65713\,
            PADIN => \N__65712\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_118_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65705\,
            DIN => \N__65704\,
            DOUT => \N__65703\,
            PACKAGEPIN => \ICE_IOR_118_wire\
        );

    \ipInertedIOPad_ICE_IOR_118_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65705\,
            PADOUT => \N__65704\,
            PADIN => \N__65703\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDO_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65696\,
            DIN => \N__65695\,
            DOUT => \N__65694\,
            PACKAGEPIN => \RTD_SDO_wire\
        );

    \ipInertedIOPad_RTD_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65696\,
            PADOUT => \N__65695\,
            PADIN => \N__65694\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65687\,
            DIN => \N__65686\,
            DOUT => \N__65685\,
            PACKAGEPIN => \IAC_OSR0_wire\
        );

    \ipInertedIOPad_IAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65687\,
            PADOUT => \N__65686\,
            PADIN => \N__65685\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__37087\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65678\,
            DIN => \N__65677\,
            DOUT => \N__65676\,
            PACKAGEPIN => \VDC_SCLK_wire\
        );

    \ipInertedIOPad_VDC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65678\,
            PADOUT => \N__65677\,
            PADIN => \N__65676\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24877\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65669\,
            DIN => \N__65668\,
            DOUT => \N__65667\,
            PACKAGEPIN => \VAC_FLT1_wire\
        );

    \ipInertedIOPad_VAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65669\,
            PADOUT => \N__65668\,
            PADIN => \N__65667\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31618\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65660\,
            DIN => \N__65659\,
            DOUT => \N__65658\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65660\,
            PADOUT => \N__65659\,
            PADIN => \N__65658\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_165_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65651\,
            DIN => \N__65650\,
            DOUT => \N__65649\,
            PACKAGEPIN => \ICE_IOR_165_wire\
        );

    \ipInertedIOPad_ICE_IOR_165_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65651\,
            PADOUT => \N__65650\,
            PADIN => \N__65649\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_147_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65642\,
            DIN => \N__65641\,
            DOUT => \N__65640\,
            PACKAGEPIN => \ICE_IOR_147_wire\
        );

    \ipInertedIOPad_ICE_IOR_147_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65642\,
            PADOUT => \N__65641\,
            PADIN => \N__65640\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_14A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65633\,
            DIN => \N__65632\,
            DOUT => \N__65631\,
            PACKAGEPIN => \ICE_IOL_14A_wire\
        );

    \ipInertedIOPad_ICE_IOL_14A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65633\,
            PADOUT => \N__65632\,
            PADIN => \N__65631\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65624\,
            DIN => \N__65623\,
            DOUT => \N__65622\,
            PACKAGEPIN => \ICE_IOL_13B_wire\
        );

    \ipInertedIOPad_ICE_IOL_13B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65624\,
            PADOUT => \N__65623\,
            PADIN => \N__65622\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_91_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65615\,
            DIN => \N__65614\,
            DOUT => \N__65613\,
            PACKAGEPIN => \ICE_IOB_91_wire\
        );

    \ipInertedIOPad_ICE_IOB_91_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65615\,
            PADOUT => \N__65614\,
            PADIN => \N__65613\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65606\,
            DIN => \N__65605\,
            DOUT => \N__65604\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65606\,
            PADOUT => \N__65605\,
            PADIN => \N__65604\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_RNG_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65597\,
            DIN => \N__65596\,
            DOUT => \N__65595\,
            PACKAGEPIN => \DDS_RNG_0_wire\
        );

    \ipInertedIOPad_DDS_RNG_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65597\,
            PADOUT => \N__65596\,
            PADIN => \N__65595\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__49897\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_RNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65588\,
            DIN => \N__65587\,
            DOUT => \N__65586\,
            PACKAGEPIN => \VDC_RNG0_wire\
        );

    \ipInertedIOPad_VDC_RNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65588\,
            PADOUT => \N__65587\,
            PADIN => \N__65586\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39892\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65579\,
            DIN => \N__65578\,
            DOUT => \N__65577\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65579\,
            PADOUT => \N__65578\,
            PADIN => \N__65577\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_152_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65570\,
            DIN => \N__65569\,
            DOUT => \N__65568\,
            PACKAGEPIN => \ICE_IOR_152_wire\
        );

    \ipInertedIOPad_ICE_IOR_152_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65570\,
            PADOUT => \N__65569\,
            PADIN => \N__65568\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65561\,
            DIN => \N__65560\,
            DOUT => \N__65559\,
            PACKAGEPIN => \ICE_IOL_12A_wire\
        );

    \ipInertedIOPad_ICE_IOL_12A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65561\,
            PADOUT => \N__65560\,
            PADIN => \N__65559\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_DRDY_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65552\,
            DIN => \N__65551\,
            DOUT => \N__65550\,
            PACKAGEPIN => \RTD_DRDY_wire\
        );

    \ipInertedIOPad_RTD_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65552\,
            PADOUT => \N__65551\,
            PADIN => \N__65550\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65543\,
            DIN => \N__65542\,
            DOUT => \N__65541\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65543\,
            PADOUT => \N__65542\,
            PADIN => \N__65541\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__35257\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_177_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65534\,
            DIN => \N__65533\,
            DOUT => \N__65532\,
            PACKAGEPIN => \ICE_IOT_177_wire\
        );

    \ipInertedIOPad_ICE_IOT_177_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65534\,
            PADOUT => \N__65533\,
            PADIN => \N__65532\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_141_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65525\,
            DIN => \N__65524\,
            DOUT => \N__65523\,
            PACKAGEPIN => \ICE_IOR_141_wire\
        );

    \ipInertedIOPad_ICE_IOR_141_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65525\,
            PADOUT => \N__65524\,
            PADIN => \N__65523\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_80_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65516\,
            DIN => \N__65515\,
            DOUT => \N__65514\,
            PACKAGEPIN => \ICE_IOB_80_wire\
        );

    \ipInertedIOPad_ICE_IOB_80_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65516\,
            PADOUT => \N__65515\,
            PADIN => \N__65514\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_102_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65507\,
            DIN => \N__65506\,
            DOUT => \N__65505\,
            PACKAGEPIN => \ICE_IOB_102_wire\
        );

    \ipInertedIOPad_ICE_IOB_102_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65507\,
            PADOUT => \N__65506\,
            PADIN => \N__65505\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65498\,
            DIN => \N__65497\,
            DOUT => \N__65496\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65498\,
            PADOUT => \N__65497\,
            PADIN => \N__65496\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65489\,
            DIN => \N__65488\,
            DOUT => \N__65487\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65489\,
            PADOUT => \N__65488\,
            PADIN => \N__65487\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__64132\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65480\,
            DIN => \N__65479\,
            DOUT => \N__65478\,
            PACKAGEPIN => \IAC_MISO_wire\
        );

    \ipInertedIOPad_IAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65480\,
            PADOUT => \N__65479\,
            PADIN => \N__65478\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65471\,
            DIN => \N__65470\,
            DOUT => \N__65469\,
            PACKAGEPIN => \VAC_OSR0_wire\
        );

    \ipInertedIOPad_VAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65471\,
            PADOUT => \N__65470\,
            PADIN => \N__65469\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__38803\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65462\,
            DIN => \N__65461\,
            DOUT => \N__65460\,
            PACKAGEPIN => \VAC_MOSI_wire\
        );

    \ipInertedIOPad_VAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65462\,
            PADOUT => \N__65461\,
            PADIN => \N__65460\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65453\,
            DIN => \N__65452\,
            DOUT => \N__65451\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65453\,
            PADOUT => \N__65452\,
            PADIN => \N__65451\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42808\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_148_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65444\,
            DIN => \N__65443\,
            DOUT => \N__65442\,
            PACKAGEPIN => \ICE_IOR_148_wire\
        );

    \ipInertedIOPad_ICE_IOR_148_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65444\,
            PADOUT => \N__65443\,
            PADIN => \N__65442\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_STAT_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65435\,
            DIN => \N__65434\,
            DOUT => \N__65433\,
            PACKAGEPIN => \STAT_COMM_wire\
        );

    \ipInertedIOPad_STAT_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65435\,
            PADOUT => \N__65434\,
            PADIN => \N__65433\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21241\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65426\,
            DIN => \N__65425\,
            DOUT => \N__65424\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65426\,
            PADOUT => \N__65425\,
            PADIN => \N__65424\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_161_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65417\,
            DIN => \N__65416\,
            DOUT => \N__65415\,
            PACKAGEPIN => \ICE_IOR_161_wire\
        );

    \ipInertedIOPad_ICE_IOR_161_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65417\,
            PADOUT => \N__65416\,
            PADIN => \N__65415\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_95_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65408\,
            DIN => \N__65407\,
            DOUT => \N__65406\,
            PACKAGEPIN => \ICE_IOB_95_wire\
        );

    \ipInertedIOPad_ICE_IOB_95_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65408\,
            PADOUT => \N__65407\,
            PADIN => \N__65406\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_82_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65399\,
            DIN => \N__65398\,
            DOUT => \N__65397\,
            PACKAGEPIN => \ICE_IOB_82_wire\
        );

    \ipInertedIOPad_ICE_IOB_82_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65399\,
            PADOUT => \N__65398\,
            PADIN => \N__65397\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_104_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65390\,
            DIN => \N__65389\,
            DOUT => \N__65388\,
            PACKAGEPIN => \ICE_IOB_104_wire\
        );

    \ipInertedIOPad_ICE_IOB_104_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65390\,
            PADOUT => \N__65389\,
            PADIN => \N__65388\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65381\,
            DIN => \N__65380\,
            DOUT => \N__65379\,
            PACKAGEPIN => \IAC_CLK_wire\
        );

    \ipInertedIOPad_IAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65381\,
            PADOUT => \N__65380\,
            PADIN => \N__65379\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26025\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65372\,
            DIN => \N__65371\,
            DOUT => \N__65370\,
            PACKAGEPIN => \DDS_CS_wire\
        );

    \ipInertedIOPad_DDS_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65372\,
            PADOUT => \N__65371\,
            PADIN => \N__65370\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__50263\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65363\,
            DIN => \N__65362\,
            DOUT => \N__65361\,
            PACKAGEPIN => \SELIRNG0_wire\
        );

    \ipInertedIOPad_SELIRNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65363\,
            PADOUT => \N__65362\,
            PADIN => \N__65361\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39943\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65354\,
            DIN => \N__65353\,
            DOUT => \N__65352\,
            PACKAGEPIN => \RTD_SDI_wire\
        );

    \ipInertedIOPad_RTD_SDI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65354\,
            PADOUT => \N__65353\,
            PADIN => \N__65352\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21280\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_221_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65345\,
            DIN => \N__65344\,
            DOUT => \N__65343\,
            PACKAGEPIN => \ICE_IOT_221_wire\
        );

    \ipInertedIOPad_ICE_IOT_221_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65345\,
            PADOUT => \N__65344\,
            PADIN => \N__65343\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_197_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65336\,
            DIN => \N__65335\,
            DOUT => \N__65334\,
            PACKAGEPIN => \ICE_IOT_197_wire\
        );

    \ipInertedIOPad_ICE_IOT_197_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65336\,
            PADOUT => \N__65335\,
            PADIN => \N__65334\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65327\,
            DIN => \N__65326\,
            DOUT => \N__65325\,
            PACKAGEPIN => \DDS_MCLK_wire\
        );

    \ipInertedIOPad_DDS_MCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65327\,
            PADOUT => \N__65326\,
            PADIN => \N__65325\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__53380\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65318\,
            DIN => \N__65317\,
            DOUT => \N__65316\,
            PACKAGEPIN => \RTD_SCLK_wire\
        );

    \ipInertedIOPad_RTD_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65318\,
            PADOUT => \N__65317\,
            PADIN => \N__65316\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21304\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65309\,
            DIN => \N__65308\,
            DOUT => \N__65307\,
            PACKAGEPIN => \RTD_CS_wire\
        );

    \ipInertedIOPad_RTD_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65309\,
            PADOUT => \N__65308\,
            PADIN => \N__65307\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22243\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_137_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65300\,
            DIN => \N__65299\,
            DOUT => \N__65298\,
            PACKAGEPIN => \ICE_IOR_137_wire\
        );

    \ipInertedIOPad_ICE_IOR_137_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65300\,
            PADOUT => \N__65299\,
            PADIN => \N__65298\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65291\,
            DIN => \N__65290\,
            DOUT => \N__65289\,
            PACKAGEPIN => \IAC_OSR1_wire\
        );

    \ipInertedIOPad_IAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65291\,
            PADOUT => \N__65290\,
            PADIN => \N__65289\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__37054\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65282\,
            DIN => \N__65281\,
            DOUT => \N__65280\,
            PACKAGEPIN => \VAC_FLT0_wire\
        );

    \ipInertedIOPad_VAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65282\,
            PADOUT => \N__65281\,
            PADIN => \N__65280\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31654\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_144_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65273\,
            DIN => \N__65272\,
            DOUT => \N__65271\,
            PACKAGEPIN => \ICE_IOR_144_wire\
        );

    \ipInertedIOPad_ICE_IOR_144_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65273\,
            PADOUT => \N__65272\,
            PADIN => \N__65271\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_128_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65264\,
            DIN => \N__65263\,
            DOUT => \N__65262\,
            PACKAGEPIN => \ICE_IOR_128_wire\
        );

    \ipInertedIOPad_ICE_IOR_128_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65264\,
            PADOUT => \N__65263\,
            PADIN => \N__65262\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65255\,
            DIN => \N__65254\,
            DOUT => \N__65253\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65255\,
            PADOUT => \N__65254\,
            PADIN => \N__65253\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65246\,
            DIN => \N__65245\,
            DOUT => \N__65244\,
            PACKAGEPIN => \IAC_SCLK_wire\
        );

    \ipInertedIOPad_IAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65246\,
            PADOUT => \N__65245\,
            PADIN => \N__65244\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27889\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65237\,
            DIN => \N__65236\,
            DOUT => \N__65235\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65237\,
            PADOUT => \N__65236\,
            PADIN => \N__65235\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \EIS_SYNCCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_139_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65228\,
            DIN => \N__65227\,
            DOUT => \N__65226\,
            PACKAGEPIN => \ICE_IOR_139_wire\
        );

    \ipInertedIOPad_ICE_IOR_139_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65228\,
            PADOUT => \N__65227\,
            PADIN => \N__65226\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65219\,
            DIN => \N__65218\,
            DOUT => \N__65217\,
            PACKAGEPIN => \ICE_IOL_4A_wire\
        );

    \ipInertedIOPad_ICE_IOL_4A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65219\,
            PADOUT => \N__65218\,
            PADIN => \N__65217\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65210\,
            DIN => \N__65209\,
            DOUT => \N__65208\,
            PACKAGEPIN => \VAC_SCLK_wire\
        );

    \ipInertedIOPad_VAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65210\,
            PADOUT => \N__65209\,
            PADIN => \N__65208\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21382\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_THERMOSTAT_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65201\,
            DIN => \N__65200\,
            DOUT => \N__65199\,
            PACKAGEPIN => \THERMOSTAT_wire\
        );

    \ipInertedIOPad_THERMOSTAT_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65201\,
            PADOUT => \N__65200\,
            PADIN => \N__65199\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \THERMOSTAT\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_164_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65192\,
            DIN => \N__65191\,
            DOUT => \N__65190\,
            PACKAGEPIN => \ICE_IOR_164_wire\
        );

    \ipInertedIOPad_ICE_IOR_164_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65192\,
            PADOUT => \N__65191\,
            PADIN => \N__65190\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_103_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65183\,
            DIN => \N__65182\,
            DOUT => \N__65181\,
            PACKAGEPIN => \ICE_IOB_103_wire\
        );

    \ipInertedIOPad_ICE_IOB_103_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65183\,
            PADOUT => \N__65182\,
            PADIN => \N__65181\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AMPV_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65174\,
            DIN => \N__65173\,
            DOUT => \N__65172\,
            PACKAGEPIN => \AMPV_POW_wire\
        );

    \ipInertedIOPad_AMPV_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65174\,
            PADOUT => \N__65173\,
            PADIN => \N__65172\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36514\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SDO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65165\,
            DIN => \N__65164\,
            DOUT => \N__65163\,
            PACKAGEPIN => \VDC_SDO_wire\
        );

    \ipInertedIOPad_VDC_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65165\,
            PADOUT => \N__65164\,
            PADIN => \N__65163\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VDC_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_174_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65156\,
            DIN => \N__65155\,
            DOUT => \N__65154\,
            PACKAGEPIN => \ICE_IOT_174_wire\
        );

    \ipInertedIOPad_ICE_IOT_174_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65156\,
            PADOUT => \N__65155\,
            PADIN => \N__65154\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_140_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65147\,
            DIN => \N__65146\,
            DOUT => \N__65145\,
            PACKAGEPIN => \ICE_IOR_140_wire\
        );

    \ipInertedIOPad_ICE_IOR_140_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65147\,
            PADOUT => \N__65146\,
            PADIN => \N__65145\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_96_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65138\,
            DIN => \N__65137\,
            DOUT => \N__65136\,
            PACKAGEPIN => \ICE_IOB_96_wire\
        );

    \ipInertedIOPad_ICE_IOB_96_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65138\,
            PADOUT => \N__65137\,
            PADIN => \N__65136\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CONT_SD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65129\,
            DIN => \N__65128\,
            DOUT => \N__65127\,
            PACKAGEPIN => \CONT_SD_wire\
        );

    \ipInertedIOPad_CONT_SD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65129\,
            PADOUT => \N__65128\,
            PADIN => \N__65127\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__52606\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AC_ADC_SYNC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65120\,
            DIN => \N__65119\,
            DOUT => \N__65118\,
            PACKAGEPIN => \AC_ADC_SYNC_wire\
        );

    \ipInertedIOPad_AC_ADC_SYNC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65120\,
            PADOUT => \N__65119\,
            PADIN => \N__65118\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23071\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65111\,
            DIN => \N__65110\,
            DOUT => \N__65109\,
            PACKAGEPIN => \SELIRNG1_wire\
        );

    \ipInertedIOPad_SELIRNG1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65111\,
            PADOUT => \N__65110\,
            PADIN => \N__65109\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__52780\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65102\,
            DIN => \N__65101\,
            DOUT => \N__65100\,
            PACKAGEPIN => \ICE_IOL_12B_wire\
        );

    \ipInertedIOPad_ICE_IOL_12B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65102\,
            PADOUT => \N__65101\,
            PADIN => \N__65100\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_160_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65093\,
            DIN => \N__65092\,
            DOUT => \N__65091\,
            PACKAGEPIN => \ICE_IOR_160_wire\
        );

    \ipInertedIOPad_ICE_IOR_160_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65093\,
            PADOUT => \N__65092\,
            PADIN => \N__65091\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_136_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65084\,
            DIN => \N__65083\,
            DOUT => \N__65082\,
            PACKAGEPIN => \ICE_IOR_136_wire\
        );

    \ipInertedIOPad_ICE_IOR_136_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65084\,
            PADOUT => \N__65083\,
            PADIN => \N__65082\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65075\,
            DIN => \N__65074\,
            DOUT => \N__65073\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65075\,
            PADOUT => \N__65074\,
            PADIN => \N__65073\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24829\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_198_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65066\,
            DIN => \N__65065\,
            DOUT => \N__65064\,
            PACKAGEPIN => \ICE_IOT_198_wire\
        );

    \ipInertedIOPad_ICE_IOT_198_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65066\,
            PADOUT => \N__65065\,
            PADIN => \N__65064\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_173_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65057\,
            DIN => \N__65056\,
            DOUT => \N__65055\,
            PACKAGEPIN => \ICE_IOT_173_wire\
        );

    \ipInertedIOPad_ICE_IOT_173_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65057\,
            PADOUT => \N__65056\,
            PADIN => \N__65055\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65048\,
            DIN => \N__65047\,
            DOUT => \N__65046\,
            PACKAGEPIN => \IAC_DRDY_wire\
        );

    \ipInertedIOPad_IAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65048\,
            PADOUT => \N__65047\,
            PADIN => \N__65046\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_178_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65039\,
            DIN => \N__65038\,
            DOUT => \N__65037\,
            PACKAGEPIN => \ICE_IOT_178_wire\
        );

    \ipInertedIOPad_ICE_IOT_178_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65039\,
            PADOUT => \N__65038\,
            PADIN => \N__65037\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_138_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65030\,
            DIN => \N__65029\,
            DOUT => \N__65028\,
            PACKAGEPIN => \ICE_IOR_138_wire\
        );

    \ipInertedIOPad_ICE_IOR_138_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65030\,
            PADOUT => \N__65029\,
            PADIN => \N__65028\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_120_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__65021\,
            DIN => \N__65020\,
            DOUT => \N__65019\,
            PACKAGEPIN => \ICE_IOR_120_wire\
        );

    \ipInertedIOPad_ICE_IOR_120_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65021\,
            PADOUT => \N__65020\,
            PADIN => \N__65019\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65012\,
            DIN => \N__65011\,
            DOUT => \N__65010\,
            PACKAGEPIN => \IAC_FLT0_wire\
        );

    \ipInertedIOPad_IAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65012\,
            PADOUT => \N__65011\,
            PADIN => \N__65010\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30574\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__65003\,
            DIN => \N__65002\,
            DOUT => \N__65001\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__65003\,
            PADOUT => \N__65002\,
            PADIN => \N__65001\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21331\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__16328\ : CascadeMux
    port map (
            O => \N__64984\,
            I => \N__64981\
        );

    \I__16327\ : InMux
    port map (
            O => \N__64981\,
            I => \N__64977\
        );

    \I__16326\ : InMux
    port map (
            O => \N__64980\,
            I => \N__64974\
        );

    \I__16325\ : LocalMux
    port map (
            O => \N__64977\,
            I => \N__64971\
        );

    \I__16324\ : LocalMux
    port map (
            O => \N__64974\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__16323\ : Odrv4
    port map (
            O => \N__64971\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__16322\ : InMux
    port map (
            O => \N__64966\,
            I => \bfn_23_6_0_\
        );

    \I__16321\ : InMux
    port map (
            O => \N__64963\,
            I => \N__64959\
        );

    \I__16320\ : InMux
    port map (
            O => \N__64962\,
            I => \N__64956\
        );

    \I__16319\ : LocalMux
    port map (
            O => \N__64959\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__16318\ : LocalMux
    port map (
            O => \N__64956\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__16317\ : InMux
    port map (
            O => \N__64951\,
            I => \ADC_VDC.genclk.n20744\
        );

    \I__16316\ : InMux
    port map (
            O => \N__64948\,
            I => \N__64944\
        );

    \I__16315\ : InMux
    port map (
            O => \N__64947\,
            I => \N__64941\
        );

    \I__16314\ : LocalMux
    port map (
            O => \N__64944\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__16313\ : LocalMux
    port map (
            O => \N__64941\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__16312\ : InMux
    port map (
            O => \N__64936\,
            I => \ADC_VDC.genclk.n20745\
        );

    \I__16311\ : InMux
    port map (
            O => \N__64933\,
            I => \N__64929\
        );

    \I__16310\ : InMux
    port map (
            O => \N__64932\,
            I => \N__64926\
        );

    \I__16309\ : LocalMux
    port map (
            O => \N__64929\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__16308\ : LocalMux
    port map (
            O => \N__64926\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__16307\ : InMux
    port map (
            O => \N__64921\,
            I => \ADC_VDC.genclk.n20746\
        );

    \I__16306\ : InMux
    port map (
            O => \N__64918\,
            I => \N__64914\
        );

    \I__16305\ : InMux
    port map (
            O => \N__64917\,
            I => \N__64911\
        );

    \I__16304\ : LocalMux
    port map (
            O => \N__64914\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__16303\ : LocalMux
    port map (
            O => \N__64911\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__16302\ : InMux
    port map (
            O => \N__64906\,
            I => \ADC_VDC.genclk.n20747\
        );

    \I__16301\ : InMux
    port map (
            O => \N__64903\,
            I => \N__64899\
        );

    \I__16300\ : InMux
    port map (
            O => \N__64902\,
            I => \N__64896\
        );

    \I__16299\ : LocalMux
    port map (
            O => \N__64899\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__16298\ : LocalMux
    port map (
            O => \N__64896\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__16297\ : InMux
    port map (
            O => \N__64891\,
            I => \ADC_VDC.genclk.n20748\
        );

    \I__16296\ : InMux
    port map (
            O => \N__64888\,
            I => \N__64884\
        );

    \I__16295\ : InMux
    port map (
            O => \N__64887\,
            I => \N__64881\
        );

    \I__16294\ : LocalMux
    port map (
            O => \N__64884\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__16293\ : LocalMux
    port map (
            O => \N__64881\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__16292\ : InMux
    port map (
            O => \N__64876\,
            I => \ADC_VDC.genclk.n20749\
        );

    \I__16291\ : SRMux
    port map (
            O => \N__64873\,
            I => \N__64870\
        );

    \I__16290\ : LocalMux
    port map (
            O => \N__64870\,
            I => \N__64865\
        );

    \I__16289\ : SRMux
    port map (
            O => \N__64869\,
            I => \N__64862\
        );

    \I__16288\ : SRMux
    port map (
            O => \N__64868\,
            I => \N__64859\
        );

    \I__16287\ : Span4Mux_v
    port map (
            O => \N__64865\,
            I => \N__64841\
        );

    \I__16286\ : LocalMux
    port map (
            O => \N__64862\,
            I => \N__64836\
        );

    \I__16285\ : LocalMux
    port map (
            O => \N__64859\,
            I => \N__64836\
        );

    \I__16284\ : SRMux
    port map (
            O => \N__64858\,
            I => \N__64833\
        );

    \I__16283\ : SRMux
    port map (
            O => \N__64857\,
            I => \N__64830\
        );

    \I__16282\ : SRMux
    port map (
            O => \N__64856\,
            I => \N__64825\
        );

    \I__16281\ : IoInMux
    port map (
            O => \N__64855\,
            I => \N__64820\
        );

    \I__16280\ : CascadeMux
    port map (
            O => \N__64854\,
            I => \N__64816\
        );

    \I__16279\ : CascadeMux
    port map (
            O => \N__64853\,
            I => \N__64812\
        );

    \I__16278\ : CascadeMux
    port map (
            O => \N__64852\,
            I => \N__64808\
        );

    \I__16277\ : CascadeMux
    port map (
            O => \N__64851\,
            I => \N__64804\
        );

    \I__16276\ : CascadeMux
    port map (
            O => \N__64850\,
            I => \N__64800\
        );

    \I__16275\ : CascadeMux
    port map (
            O => \N__64849\,
            I => \N__64796\
        );

    \I__16274\ : CascadeMux
    port map (
            O => \N__64848\,
            I => \N__64792\
        );

    \I__16273\ : CascadeMux
    port map (
            O => \N__64847\,
            I => \N__64789\
        );

    \I__16272\ : CascadeMux
    port map (
            O => \N__64846\,
            I => \N__64785\
        );

    \I__16271\ : CascadeMux
    port map (
            O => \N__64845\,
            I => \N__64781\
        );

    \I__16270\ : CascadeMux
    port map (
            O => \N__64844\,
            I => \N__64777\
        );

    \I__16269\ : Span4Mux_v
    port map (
            O => \N__64841\,
            I => \N__64774\
        );

    \I__16268\ : Span4Mux_v
    port map (
            O => \N__64836\,
            I => \N__64767\
        );

    \I__16267\ : LocalMux
    port map (
            O => \N__64833\,
            I => \N__64767\
        );

    \I__16266\ : LocalMux
    port map (
            O => \N__64830\,
            I => \N__64767\
        );

    \I__16265\ : SRMux
    port map (
            O => \N__64829\,
            I => \N__64764\
        );

    \I__16264\ : SRMux
    port map (
            O => \N__64828\,
            I => \N__64761\
        );

    \I__16263\ : LocalMux
    port map (
            O => \N__64825\,
            I => \N__64758\
        );

    \I__16262\ : SRMux
    port map (
            O => \N__64824\,
            I => \N__64755\
        );

    \I__16261\ : SRMux
    port map (
            O => \N__64823\,
            I => \N__64752\
        );

    \I__16260\ : LocalMux
    port map (
            O => \N__64820\,
            I => \N__64749\
        );

    \I__16259\ : InMux
    port map (
            O => \N__64819\,
            I => \N__64734\
        );

    \I__16258\ : InMux
    port map (
            O => \N__64816\,
            I => \N__64734\
        );

    \I__16257\ : InMux
    port map (
            O => \N__64815\,
            I => \N__64734\
        );

    \I__16256\ : InMux
    port map (
            O => \N__64812\,
            I => \N__64734\
        );

    \I__16255\ : InMux
    port map (
            O => \N__64811\,
            I => \N__64734\
        );

    \I__16254\ : InMux
    port map (
            O => \N__64808\,
            I => \N__64734\
        );

    \I__16253\ : InMux
    port map (
            O => \N__64807\,
            I => \N__64734\
        );

    \I__16252\ : InMux
    port map (
            O => \N__64804\,
            I => \N__64712\
        );

    \I__16251\ : InMux
    port map (
            O => \N__64803\,
            I => \N__64712\
        );

    \I__16250\ : InMux
    port map (
            O => \N__64800\,
            I => \N__64712\
        );

    \I__16249\ : InMux
    port map (
            O => \N__64799\,
            I => \N__64712\
        );

    \I__16248\ : InMux
    port map (
            O => \N__64796\,
            I => \N__64712\
        );

    \I__16247\ : InMux
    port map (
            O => \N__64795\,
            I => \N__64712\
        );

    \I__16246\ : InMux
    port map (
            O => \N__64792\,
            I => \N__64712\
        );

    \I__16245\ : InMux
    port map (
            O => \N__64789\,
            I => \N__64697\
        );

    \I__16244\ : InMux
    port map (
            O => \N__64788\,
            I => \N__64697\
        );

    \I__16243\ : InMux
    port map (
            O => \N__64785\,
            I => \N__64697\
        );

    \I__16242\ : InMux
    port map (
            O => \N__64784\,
            I => \N__64697\
        );

    \I__16241\ : InMux
    port map (
            O => \N__64781\,
            I => \N__64697\
        );

    \I__16240\ : InMux
    port map (
            O => \N__64780\,
            I => \N__64697\
        );

    \I__16239\ : InMux
    port map (
            O => \N__64777\,
            I => \N__64697\
        );

    \I__16238\ : Span4Mux_v
    port map (
            O => \N__64774\,
            I => \N__64684\
        );

    \I__16237\ : Span4Mux_v
    port map (
            O => \N__64767\,
            I => \N__64684\
        );

    \I__16236\ : LocalMux
    port map (
            O => \N__64764\,
            I => \N__64684\
        );

    \I__16235\ : LocalMux
    port map (
            O => \N__64761\,
            I => \N__64684\
        );

    \I__16234\ : Span4Mux_v
    port map (
            O => \N__64758\,
            I => \N__64677\
        );

    \I__16233\ : LocalMux
    port map (
            O => \N__64755\,
            I => \N__64677\
        );

    \I__16232\ : LocalMux
    port map (
            O => \N__64752\,
            I => \N__64677\
        );

    \I__16231\ : Span4Mux_s3_v
    port map (
            O => \N__64749\,
            I => \N__64673\
        );

    \I__16230\ : LocalMux
    port map (
            O => \N__64734\,
            I => \N__64670\
        );

    \I__16229\ : CascadeMux
    port map (
            O => \N__64733\,
            I => \N__64667\
        );

    \I__16228\ : CascadeMux
    port map (
            O => \N__64732\,
            I => \N__64663\
        );

    \I__16227\ : CascadeMux
    port map (
            O => \N__64731\,
            I => \N__64660\
        );

    \I__16226\ : CascadeMux
    port map (
            O => \N__64730\,
            I => \N__64657\
        );

    \I__16225\ : CascadeMux
    port map (
            O => \N__64729\,
            I => \N__64654\
        );

    \I__16224\ : CascadeMux
    port map (
            O => \N__64728\,
            I => \N__64651\
        );

    \I__16223\ : CascadeMux
    port map (
            O => \N__64727\,
            I => \N__64648\
        );

    \I__16222\ : LocalMux
    port map (
            O => \N__64712\,
            I => \N__64645\
        );

    \I__16221\ : LocalMux
    port map (
            O => \N__64697\,
            I => \N__64642\
        );

    \I__16220\ : CascadeMux
    port map (
            O => \N__64696\,
            I => \N__64638\
        );

    \I__16219\ : CascadeMux
    port map (
            O => \N__64695\,
            I => \N__64634\
        );

    \I__16218\ : CascadeMux
    port map (
            O => \N__64694\,
            I => \N__64630\
        );

    \I__16217\ : CascadeMux
    port map (
            O => \N__64693\,
            I => \N__64626\
        );

    \I__16216\ : Span4Mux_v
    port map (
            O => \N__64684\,
            I => \N__64621\
        );

    \I__16215\ : Span4Mux_v
    port map (
            O => \N__64677\,
            I => \N__64621\
        );

    \I__16214\ : InMux
    port map (
            O => \N__64676\,
            I => \N__64618\
        );

    \I__16213\ : Span4Mux_v
    port map (
            O => \N__64673\,
            I => \N__64613\
        );

    \I__16212\ : Span4Mux_h
    port map (
            O => \N__64670\,
            I => \N__64610\
        );

    \I__16211\ : InMux
    port map (
            O => \N__64667\,
            I => \N__64601\
        );

    \I__16210\ : InMux
    port map (
            O => \N__64666\,
            I => \N__64601\
        );

    \I__16209\ : InMux
    port map (
            O => \N__64663\,
            I => \N__64601\
        );

    \I__16208\ : InMux
    port map (
            O => \N__64660\,
            I => \N__64601\
        );

    \I__16207\ : InMux
    port map (
            O => \N__64657\,
            I => \N__64592\
        );

    \I__16206\ : InMux
    port map (
            O => \N__64654\,
            I => \N__64592\
        );

    \I__16205\ : InMux
    port map (
            O => \N__64651\,
            I => \N__64592\
        );

    \I__16204\ : InMux
    port map (
            O => \N__64648\,
            I => \N__64592\
        );

    \I__16203\ : Span4Mux_v
    port map (
            O => \N__64645\,
            I => \N__64587\
        );

    \I__16202\ : Span4Mux_v
    port map (
            O => \N__64642\,
            I => \N__64587\
        );

    \I__16201\ : InMux
    port map (
            O => \N__64641\,
            I => \N__64570\
        );

    \I__16200\ : InMux
    port map (
            O => \N__64638\,
            I => \N__64570\
        );

    \I__16199\ : InMux
    port map (
            O => \N__64637\,
            I => \N__64570\
        );

    \I__16198\ : InMux
    port map (
            O => \N__64634\,
            I => \N__64570\
        );

    \I__16197\ : InMux
    port map (
            O => \N__64633\,
            I => \N__64570\
        );

    \I__16196\ : InMux
    port map (
            O => \N__64630\,
            I => \N__64570\
        );

    \I__16195\ : InMux
    port map (
            O => \N__64629\,
            I => \N__64570\
        );

    \I__16194\ : InMux
    port map (
            O => \N__64626\,
            I => \N__64570\
        );

    \I__16193\ : Span4Mux_h
    port map (
            O => \N__64621\,
            I => \N__64567\
        );

    \I__16192\ : LocalMux
    port map (
            O => \N__64618\,
            I => \N__64564\
        );

    \I__16191\ : SRMux
    port map (
            O => \N__64617\,
            I => \N__64561\
        );

    \I__16190\ : SRMux
    port map (
            O => \N__64616\,
            I => \N__64558\
        );

    \I__16189\ : Span4Mux_v
    port map (
            O => \N__64613\,
            I => \N__64554\
        );

    \I__16188\ : Sp12to4
    port map (
            O => \N__64610\,
            I => \N__64551\
        );

    \I__16187\ : LocalMux
    port map (
            O => \N__64601\,
            I => \N__64542\
        );

    \I__16186\ : LocalMux
    port map (
            O => \N__64592\,
            I => \N__64542\
        );

    \I__16185\ : Sp12to4
    port map (
            O => \N__64587\,
            I => \N__64542\
        );

    \I__16184\ : LocalMux
    port map (
            O => \N__64570\,
            I => \N__64542\
        );

    \I__16183\ : Span4Mux_h
    port map (
            O => \N__64567\,
            I => \N__64537\
        );

    \I__16182\ : Span4Mux_v
    port map (
            O => \N__64564\,
            I => \N__64537\
        );

    \I__16181\ : LocalMux
    port map (
            O => \N__64561\,
            I => \N__64534\
        );

    \I__16180\ : LocalMux
    port map (
            O => \N__64558\,
            I => \N__64531\
        );

    \I__16179\ : InMux
    port map (
            O => \N__64557\,
            I => \N__64528\
        );

    \I__16178\ : Sp12to4
    port map (
            O => \N__64554\,
            I => \N__64521\
        );

    \I__16177\ : Span12Mux_v
    port map (
            O => \N__64551\,
            I => \N__64521\
        );

    \I__16176\ : Span12Mux_h
    port map (
            O => \N__64542\,
            I => \N__64521\
        );

    \I__16175\ : Span4Mux_h
    port map (
            O => \N__64537\,
            I => \N__64518\
        );

    \I__16174\ : Span4Mux_v
    port map (
            O => \N__64534\,
            I => \N__64513\
        );

    \I__16173\ : Span4Mux_v
    port map (
            O => \N__64531\,
            I => \N__64513\
        );

    \I__16172\ : LocalMux
    port map (
            O => \N__64528\,
            I => \N__64510\
        );

    \I__16171\ : Odrv12
    port map (
            O => \N__64521\,
            I => \CONSTANT_ONE_NET\
        );

    \I__16170\ : Odrv4
    port map (
            O => \N__64518\,
            I => \CONSTANT_ONE_NET\
        );

    \I__16169\ : Odrv4
    port map (
            O => \N__64513\,
            I => \CONSTANT_ONE_NET\
        );

    \I__16168\ : Odrv4
    port map (
            O => \N__64510\,
            I => \CONSTANT_ONE_NET\
        );

    \I__16167\ : InMux
    port map (
            O => \N__64501\,
            I => \ADC_VDC.genclk.n20750\
        );

    \I__16166\ : CascadeMux
    port map (
            O => \N__64498\,
            I => \N__64494\
        );

    \I__16165\ : InMux
    port map (
            O => \N__64497\,
            I => \N__64491\
        );

    \I__16164\ : InMux
    port map (
            O => \N__64494\,
            I => \N__64488\
        );

    \I__16163\ : LocalMux
    port map (
            O => \N__64491\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__16162\ : LocalMux
    port map (
            O => \N__64488\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__16161\ : CEMux
    port map (
            O => \N__64483\,
            I => \N__64480\
        );

    \I__16160\ : LocalMux
    port map (
            O => \N__64480\,
            I => \N__64476\
        );

    \I__16159\ : CEMux
    port map (
            O => \N__64479\,
            I => \N__64473\
        );

    \I__16158\ : Span4Mux_v
    port map (
            O => \N__64476\,
            I => \N__64470\
        );

    \I__16157\ : LocalMux
    port map (
            O => \N__64473\,
            I => \N__64467\
        );

    \I__16156\ : Span4Mux_h
    port map (
            O => \N__64470\,
            I => \N__64462\
        );

    \I__16155\ : Span4Mux_h
    port map (
            O => \N__64467\,
            I => \N__64462\
        );

    \I__16154\ : Odrv4
    port map (
            O => \N__64462\,
            I => \ADC_VDC.genclk.n12361\
        );

    \I__16153\ : SRMux
    port map (
            O => \N__64459\,
            I => \N__64454\
        );

    \I__16152\ : SRMux
    port map (
            O => \N__64458\,
            I => \N__64451\
        );

    \I__16151\ : SRMux
    port map (
            O => \N__64457\,
            I => \N__64448\
        );

    \I__16150\ : LocalMux
    port map (
            O => \N__64454\,
            I => \N__64444\
        );

    \I__16149\ : LocalMux
    port map (
            O => \N__64451\,
            I => \N__64441\
        );

    \I__16148\ : LocalMux
    port map (
            O => \N__64448\,
            I => \N__64438\
        );

    \I__16147\ : SRMux
    port map (
            O => \N__64447\,
            I => \N__64435\
        );

    \I__16146\ : Span4Mux_h
    port map (
            O => \N__64444\,
            I => \N__64432\
        );

    \I__16145\ : Span4Mux_h
    port map (
            O => \N__64441\,
            I => \N__64427\
        );

    \I__16144\ : Span4Mux_h
    port map (
            O => \N__64438\,
            I => \N__64427\
        );

    \I__16143\ : LocalMux
    port map (
            O => \N__64435\,
            I => \N__64424\
        );

    \I__16142\ : Odrv4
    port map (
            O => \N__64432\,
            I => \ADC_VDC.genclk.n15418\
        );

    \I__16141\ : Odrv4
    port map (
            O => \N__64427\,
            I => \ADC_VDC.genclk.n15418\
        );

    \I__16140\ : Odrv4
    port map (
            O => \N__64424\,
            I => \ADC_VDC.genclk.n15418\
        );

    \I__16139\ : SRMux
    port map (
            O => \N__64417\,
            I => \N__64413\
        );

    \I__16138\ : SRMux
    port map (
            O => \N__64416\,
            I => \N__64410\
        );

    \I__16137\ : LocalMux
    port map (
            O => \N__64413\,
            I => \N__64407\
        );

    \I__16136\ : LocalMux
    port map (
            O => \N__64410\,
            I => \N__64404\
        );

    \I__16135\ : Span4Mux_h
    port map (
            O => \N__64407\,
            I => \N__64401\
        );

    \I__16134\ : Span4Mux_h
    port map (
            O => \N__64404\,
            I => \N__64398\
        );

    \I__16133\ : Odrv4
    port map (
            O => \N__64401\,
            I => n15482
        );

    \I__16132\ : Odrv4
    port map (
            O => \N__64398\,
            I => n15482
        );

    \I__16131\ : InMux
    port map (
            O => \N__64393\,
            I => \N__64389\
        );

    \I__16130\ : InMux
    port map (
            O => \N__64392\,
            I => \N__64386\
        );

    \I__16129\ : LocalMux
    port map (
            O => \N__64389\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__16128\ : LocalMux
    port map (
            O => \N__64386\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__16127\ : InMux
    port map (
            O => \N__64381\,
            I => \bfn_23_5_0_\
        );

    \I__16126\ : InMux
    port map (
            O => \N__64378\,
            I => \N__64374\
        );

    \I__16125\ : InMux
    port map (
            O => \N__64377\,
            I => \N__64371\
        );

    \I__16124\ : LocalMux
    port map (
            O => \N__64374\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__16123\ : LocalMux
    port map (
            O => \N__64371\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__16122\ : InMux
    port map (
            O => \N__64366\,
            I => \ADC_VDC.genclk.n20736\
        );

    \I__16121\ : CascadeMux
    port map (
            O => \N__64363\,
            I => \N__64360\
        );

    \I__16120\ : InMux
    port map (
            O => \N__64360\,
            I => \N__64356\
        );

    \I__16119\ : InMux
    port map (
            O => \N__64359\,
            I => \N__64353\
        );

    \I__16118\ : LocalMux
    port map (
            O => \N__64356\,
            I => \N__64348\
        );

    \I__16117\ : LocalMux
    port map (
            O => \N__64353\,
            I => \N__64348\
        );

    \I__16116\ : Odrv4
    port map (
            O => \N__64348\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__16115\ : InMux
    port map (
            O => \N__64345\,
            I => \ADC_VDC.genclk.n20737\
        );

    \I__16114\ : InMux
    port map (
            O => \N__64342\,
            I => \N__64338\
        );

    \I__16113\ : InMux
    port map (
            O => \N__64341\,
            I => \N__64335\
        );

    \I__16112\ : LocalMux
    port map (
            O => \N__64338\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__16111\ : LocalMux
    port map (
            O => \N__64335\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__16110\ : InMux
    port map (
            O => \N__64330\,
            I => \ADC_VDC.genclk.n20738\
        );

    \I__16109\ : CascadeMux
    port map (
            O => \N__64327\,
            I => \N__64323\
        );

    \I__16108\ : CascadeMux
    port map (
            O => \N__64326\,
            I => \N__64320\
        );

    \I__16107\ : InMux
    port map (
            O => \N__64323\,
            I => \N__64317\
        );

    \I__16106\ : InMux
    port map (
            O => \N__64320\,
            I => \N__64314\
        );

    \I__16105\ : LocalMux
    port map (
            O => \N__64317\,
            I => \N__64311\
        );

    \I__16104\ : LocalMux
    port map (
            O => \N__64314\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__16103\ : Odrv4
    port map (
            O => \N__64311\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__16102\ : InMux
    port map (
            O => \N__64306\,
            I => \ADC_VDC.genclk.n20739\
        );

    \I__16101\ : InMux
    port map (
            O => \N__64303\,
            I => \N__64299\
        );

    \I__16100\ : InMux
    port map (
            O => \N__64302\,
            I => \N__64296\
        );

    \I__16099\ : LocalMux
    port map (
            O => \N__64299\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__16098\ : LocalMux
    port map (
            O => \N__64296\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__16097\ : InMux
    port map (
            O => \N__64291\,
            I => \ADC_VDC.genclk.n20740\
        );

    \I__16096\ : CascadeMux
    port map (
            O => \N__64288\,
            I => \N__64285\
        );

    \I__16095\ : InMux
    port map (
            O => \N__64285\,
            I => \N__64281\
        );

    \I__16094\ : InMux
    port map (
            O => \N__64284\,
            I => \N__64278\
        );

    \I__16093\ : LocalMux
    port map (
            O => \N__64281\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__16092\ : LocalMux
    port map (
            O => \N__64278\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__16091\ : InMux
    port map (
            O => \N__64273\,
            I => \ADC_VDC.genclk.n20741\
        );

    \I__16090\ : CascadeMux
    port map (
            O => \N__64270\,
            I => \N__64266\
        );

    \I__16089\ : InMux
    port map (
            O => \N__64269\,
            I => \N__64263\
        );

    \I__16088\ : InMux
    port map (
            O => \N__64266\,
            I => \N__64260\
        );

    \I__16087\ : LocalMux
    port map (
            O => \N__64263\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__16086\ : LocalMux
    port map (
            O => \N__64260\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__16085\ : InMux
    port map (
            O => \N__64255\,
            I => \ADC_VDC.genclk.n20742\
        );

    \I__16084\ : InMux
    port map (
            O => \N__64252\,
            I => \N__64249\
        );

    \I__16083\ : LocalMux
    port map (
            O => \N__64249\,
            I => \ADC_VDC.genclk.n26\
        );

    \I__16082\ : CascadeMux
    port map (
            O => \N__64246\,
            I => \ADC_VDC.genclk.n22305_cascade_\
        );

    \I__16081\ : InMux
    port map (
            O => \N__64243\,
            I => \N__64240\
        );

    \I__16080\ : LocalMux
    port map (
            O => \N__64240\,
            I => \ADC_VDC.genclk.n27\
        );

    \I__16079\ : InMux
    port map (
            O => \N__64237\,
            I => \N__64234\
        );

    \I__16078\ : LocalMux
    port map (
            O => \N__64234\,
            I => \N__64231\
        );

    \I__16077\ : Odrv4
    port map (
            O => \N__64231\,
            I => \ADC_VDC.genclk.n22303\
        );

    \I__16076\ : InMux
    port map (
            O => \N__64228\,
            I => \N__64224\
        );

    \I__16075\ : InMux
    port map (
            O => \N__64227\,
            I => \N__64221\
        );

    \I__16074\ : LocalMux
    port map (
            O => \N__64224\,
            I => \N__64211\
        );

    \I__16073\ : LocalMux
    port map (
            O => \N__64221\,
            I => \N__64211\
        );

    \I__16072\ : InMux
    port map (
            O => \N__64220\,
            I => \N__64206\
        );

    \I__16071\ : InMux
    port map (
            O => \N__64219\,
            I => \N__64206\
        );

    \I__16070\ : InMux
    port map (
            O => \N__64218\,
            I => \N__64203\
        );

    \I__16069\ : InMux
    port map (
            O => \N__64217\,
            I => \N__64198\
        );

    \I__16068\ : InMux
    port map (
            O => \N__64216\,
            I => \N__64198\
        );

    \I__16067\ : Odrv12
    port map (
            O => \N__64211\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__16066\ : LocalMux
    port map (
            O => \N__64206\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__16065\ : LocalMux
    port map (
            O => \N__64203\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__16064\ : LocalMux
    port map (
            O => \N__64198\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__16063\ : CascadeMux
    port map (
            O => \N__64189\,
            I => \ADC_VDC.genclk.n22303_cascade_\
        );

    \I__16062\ : InMux
    port map (
            O => \N__64186\,
            I => \N__64183\
        );

    \I__16061\ : LocalMux
    port map (
            O => \N__64183\,
            I => \N__64180\
        );

    \I__16060\ : Span4Mux_v
    port map (
            O => \N__64180\,
            I => \N__64176\
        );

    \I__16059\ : InMux
    port map (
            O => \N__64179\,
            I => \N__64173\
        );

    \I__16058\ : Odrv4
    port map (
            O => \N__64176\,
            I => \ADC_VDC.genclk.n22302\
        );

    \I__16057\ : LocalMux
    port map (
            O => \N__64173\,
            I => \ADC_VDC.genclk.n22302\
        );

    \I__16056\ : CascadeMux
    port map (
            O => \N__64168\,
            I => \N__64164\
        );

    \I__16055\ : InMux
    port map (
            O => \N__64167\,
            I => \N__64154\
        );

    \I__16054\ : InMux
    port map (
            O => \N__64164\,
            I => \N__64154\
        );

    \I__16053\ : InMux
    port map (
            O => \N__64163\,
            I => \N__64154\
        );

    \I__16052\ : InMux
    port map (
            O => \N__64162\,
            I => \N__64151\
        );

    \I__16051\ : InMux
    port map (
            O => \N__64161\,
            I => \N__64148\
        );

    \I__16050\ : LocalMux
    port map (
            O => \N__64154\,
            I => \N__64143\
        );

    \I__16049\ : LocalMux
    port map (
            O => \N__64151\,
            I => \N__64143\
        );

    \I__16048\ : LocalMux
    port map (
            O => \N__64148\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__16047\ : Odrv4
    port map (
            O => \N__64143\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__16046\ : InMux
    port map (
            O => \N__64138\,
            I => \N__64135\
        );

    \I__16045\ : LocalMux
    port map (
            O => \N__64135\,
            I => \ADC_VDC.genclk.n28\
        );

    \I__16044\ : IoInMux
    port map (
            O => \N__64132\,
            I => \N__64129\
        );

    \I__16043\ : LocalMux
    port map (
            O => \N__64129\,
            I => \N__64126\
        );

    \I__16042\ : IoSpan4Mux
    port map (
            O => \N__64126\,
            I => \N__64123\
        );

    \I__16041\ : IoSpan4Mux
    port map (
            O => \N__64123\,
            I => \N__64120\
        );

    \I__16040\ : IoSpan4Mux
    port map (
            O => \N__64120\,
            I => \N__64117\
        );

    \I__16039\ : Span4Mux_s3_h
    port map (
            O => \N__64117\,
            I => \N__64114\
        );

    \I__16038\ : Odrv4
    port map (
            O => \N__64114\,
            I => \ICE_GPMI_0\
        );

    \I__16037\ : InMux
    port map (
            O => \N__64111\,
            I => \N__64102\
        );

    \I__16036\ : InMux
    port map (
            O => \N__64110\,
            I => \N__64102\
        );

    \I__16035\ : InMux
    port map (
            O => \N__64109\,
            I => \N__64102\
        );

    \I__16034\ : LocalMux
    port map (
            O => \N__64102\,
            I => \N__64098\
        );

    \I__16033\ : CascadeMux
    port map (
            O => \N__64101\,
            I => \N__64092\
        );

    \I__16032\ : Span4Mux_v
    port map (
            O => \N__64098\,
            I => \N__64085\
        );

    \I__16031\ : InMux
    port map (
            O => \N__64097\,
            I => \N__64080\
        );

    \I__16030\ : InMux
    port map (
            O => \N__64096\,
            I => \N__64080\
        );

    \I__16029\ : InMux
    port map (
            O => \N__64095\,
            I => \N__64067\
        );

    \I__16028\ : InMux
    port map (
            O => \N__64092\,
            I => \N__64067\
        );

    \I__16027\ : InMux
    port map (
            O => \N__64091\,
            I => \N__64067\
        );

    \I__16026\ : InMux
    port map (
            O => \N__64090\,
            I => \N__64067\
        );

    \I__16025\ : InMux
    port map (
            O => \N__64089\,
            I => \N__64062\
        );

    \I__16024\ : InMux
    port map (
            O => \N__64088\,
            I => \N__64059\
        );

    \I__16023\ : Span4Mux_h
    port map (
            O => \N__64085\,
            I => \N__64054\
        );

    \I__16022\ : LocalMux
    port map (
            O => \N__64080\,
            I => \N__64054\
        );

    \I__16021\ : InMux
    port map (
            O => \N__64079\,
            I => \N__64051\
        );

    \I__16020\ : InMux
    port map (
            O => \N__64078\,
            I => \N__64041\
        );

    \I__16019\ : InMux
    port map (
            O => \N__64077\,
            I => \N__64041\
        );

    \I__16018\ : InMux
    port map (
            O => \N__64076\,
            I => \N__64041\
        );

    \I__16017\ : LocalMux
    port map (
            O => \N__64067\,
            I => \N__64038\
        );

    \I__16016\ : CascadeMux
    port map (
            O => \N__64066\,
            I => \N__64035\
        );

    \I__16015\ : InMux
    port map (
            O => \N__64065\,
            I => \N__64026\
        );

    \I__16014\ : LocalMux
    port map (
            O => \N__64062\,
            I => \N__64017\
        );

    \I__16013\ : LocalMux
    port map (
            O => \N__64059\,
            I => \N__64017\
        );

    \I__16012\ : Span4Mux_v
    port map (
            O => \N__64054\,
            I => \N__64012\
        );

    \I__16011\ : LocalMux
    port map (
            O => \N__64051\,
            I => \N__64012\
        );

    \I__16010\ : CascadeMux
    port map (
            O => \N__64050\,
            I => \N__64008\
        );

    \I__16009\ : InMux
    port map (
            O => \N__64049\,
            I => \N__64001\
        );

    \I__16008\ : InMux
    port map (
            O => \N__64048\,
            I => \N__64001\
        );

    \I__16007\ : LocalMux
    port map (
            O => \N__64041\,
            I => \N__63998\
        );

    \I__16006\ : Span4Mux_v
    port map (
            O => \N__64038\,
            I => \N__63995\
        );

    \I__16005\ : InMux
    port map (
            O => \N__64035\,
            I => \N__63980\
        );

    \I__16004\ : InMux
    port map (
            O => \N__64034\,
            I => \N__63980\
        );

    \I__16003\ : InMux
    port map (
            O => \N__64033\,
            I => \N__63973\
        );

    \I__16002\ : InMux
    port map (
            O => \N__64032\,
            I => \N__63973\
        );

    \I__16001\ : InMux
    port map (
            O => \N__64031\,
            I => \N__63973\
        );

    \I__16000\ : InMux
    port map (
            O => \N__64030\,
            I => \N__63970\
        );

    \I__15999\ : CascadeMux
    port map (
            O => \N__64029\,
            I => \N__63967\
        );

    \I__15998\ : LocalMux
    port map (
            O => \N__64026\,
            I => \N__63963\
        );

    \I__15997\ : InMux
    port map (
            O => \N__64025\,
            I => \N__63960\
        );

    \I__15996\ : InMux
    port map (
            O => \N__64024\,
            I => \N__63956\
        );

    \I__15995\ : InMux
    port map (
            O => \N__64023\,
            I => \N__63951\
        );

    \I__15994\ : InMux
    port map (
            O => \N__64022\,
            I => \N__63951\
        );

    \I__15993\ : Span4Mux_v
    port map (
            O => \N__64017\,
            I => \N__63946\
        );

    \I__15992\ : Span4Mux_v
    port map (
            O => \N__64012\,
            I => \N__63946\
        );

    \I__15991\ : InMux
    port map (
            O => \N__64011\,
            I => \N__63941\
        );

    \I__15990\ : InMux
    port map (
            O => \N__64008\,
            I => \N__63941\
        );

    \I__15989\ : InMux
    port map (
            O => \N__64007\,
            I => \N__63936\
        );

    \I__15988\ : InMux
    port map (
            O => \N__64006\,
            I => \N__63936\
        );

    \I__15987\ : LocalMux
    port map (
            O => \N__64001\,
            I => \N__63931\
        );

    \I__15986\ : Span4Mux_h
    port map (
            O => \N__63998\,
            I => \N__63931\
        );

    \I__15985\ : Span4Mux_h
    port map (
            O => \N__63995\,
            I => \N__63928\
        );

    \I__15984\ : InMux
    port map (
            O => \N__63994\,
            I => \N__63923\
        );

    \I__15983\ : InMux
    port map (
            O => \N__63993\,
            I => \N__63923\
        );

    \I__15982\ : InMux
    port map (
            O => \N__63992\,
            I => \N__63920\
        );

    \I__15981\ : InMux
    port map (
            O => \N__63991\,
            I => \N__63911\
        );

    \I__15980\ : InMux
    port map (
            O => \N__63990\,
            I => \N__63911\
        );

    \I__15979\ : InMux
    port map (
            O => \N__63989\,
            I => \N__63911\
        );

    \I__15978\ : InMux
    port map (
            O => \N__63988\,
            I => \N__63911\
        );

    \I__15977\ : CascadeMux
    port map (
            O => \N__63987\,
            I => \N__63905\
        );

    \I__15976\ : CascadeMux
    port map (
            O => \N__63986\,
            I => \N__63902\
        );

    \I__15975\ : InMux
    port map (
            O => \N__63985\,
            I => \N__63899\
        );

    \I__15974\ : LocalMux
    port map (
            O => \N__63980\,
            I => \N__63896\
        );

    \I__15973\ : LocalMux
    port map (
            O => \N__63973\,
            I => \N__63893\
        );

    \I__15972\ : LocalMux
    port map (
            O => \N__63970\,
            I => \N__63890\
        );

    \I__15971\ : InMux
    port map (
            O => \N__63967\,
            I => \N__63885\
        );

    \I__15970\ : InMux
    port map (
            O => \N__63966\,
            I => \N__63882\
        );

    \I__15969\ : Span4Mux_h
    port map (
            O => \N__63963\,
            I => \N__63879\
        );

    \I__15968\ : LocalMux
    port map (
            O => \N__63960\,
            I => \N__63876\
        );

    \I__15967\ : InMux
    port map (
            O => \N__63959\,
            I => \N__63873\
        );

    \I__15966\ : LocalMux
    port map (
            O => \N__63956\,
            I => \N__63868\
        );

    \I__15965\ : LocalMux
    port map (
            O => \N__63951\,
            I => \N__63868\
        );

    \I__15964\ : Span4Mux_h
    port map (
            O => \N__63946\,
            I => \N__63865\
        );

    \I__15963\ : LocalMux
    port map (
            O => \N__63941\,
            I => \N__63860\
        );

    \I__15962\ : LocalMux
    port map (
            O => \N__63936\,
            I => \N__63860\
        );

    \I__15961\ : Span4Mux_v
    port map (
            O => \N__63931\,
            I => \N__63853\
        );

    \I__15960\ : Span4Mux_v
    port map (
            O => \N__63928\,
            I => \N__63853\
        );

    \I__15959\ : LocalMux
    port map (
            O => \N__63923\,
            I => \N__63853\
        );

    \I__15958\ : LocalMux
    port map (
            O => \N__63920\,
            I => \N__63848\
        );

    \I__15957\ : LocalMux
    port map (
            O => \N__63911\,
            I => \N__63848\
        );

    \I__15956\ : InMux
    port map (
            O => \N__63910\,
            I => \N__63845\
        );

    \I__15955\ : InMux
    port map (
            O => \N__63909\,
            I => \N__63836\
        );

    \I__15954\ : InMux
    port map (
            O => \N__63908\,
            I => \N__63836\
        );

    \I__15953\ : InMux
    port map (
            O => \N__63905\,
            I => \N__63836\
        );

    \I__15952\ : InMux
    port map (
            O => \N__63902\,
            I => \N__63836\
        );

    \I__15951\ : LocalMux
    port map (
            O => \N__63899\,
            I => \N__63827\
        );

    \I__15950\ : Span4Mux_v
    port map (
            O => \N__63896\,
            I => \N__63827\
        );

    \I__15949\ : Span4Mux_v
    port map (
            O => \N__63893\,
            I => \N__63827\
        );

    \I__15948\ : Span4Mux_v
    port map (
            O => \N__63890\,
            I => \N__63827\
        );

    \I__15947\ : InMux
    port map (
            O => \N__63889\,
            I => \N__63822\
        );

    \I__15946\ : InMux
    port map (
            O => \N__63888\,
            I => \N__63822\
        );

    \I__15945\ : LocalMux
    port map (
            O => \N__63885\,
            I => \N__63815\
        );

    \I__15944\ : LocalMux
    port map (
            O => \N__63882\,
            I => \N__63815\
        );

    \I__15943\ : Span4Mux_h
    port map (
            O => \N__63879\,
            I => \N__63815\
        );

    \I__15942\ : Span4Mux_v
    port map (
            O => \N__63876\,
            I => \N__63802\
        );

    \I__15941\ : LocalMux
    port map (
            O => \N__63873\,
            I => \N__63802\
        );

    \I__15940\ : Span4Mux_h
    port map (
            O => \N__63868\,
            I => \N__63802\
        );

    \I__15939\ : Span4Mux_h
    port map (
            O => \N__63865\,
            I => \N__63802\
        );

    \I__15938\ : Span4Mux_v
    port map (
            O => \N__63860\,
            I => \N__63802\
        );

    \I__15937\ : Span4Mux_v
    port map (
            O => \N__63853\,
            I => \N__63802\
        );

    \I__15936\ : Span12Mux_v
    port map (
            O => \N__63848\,
            I => \N__63799\
        );

    \I__15935\ : LocalMux
    port map (
            O => \N__63845\,
            I => comm_state_2
        );

    \I__15934\ : LocalMux
    port map (
            O => \N__63836\,
            I => comm_state_2
        );

    \I__15933\ : Odrv4
    port map (
            O => \N__63827\,
            I => comm_state_2
        );

    \I__15932\ : LocalMux
    port map (
            O => \N__63822\,
            I => comm_state_2
        );

    \I__15931\ : Odrv4
    port map (
            O => \N__63815\,
            I => comm_state_2
        );

    \I__15930\ : Odrv4
    port map (
            O => \N__63802\,
            I => comm_state_2
        );

    \I__15929\ : Odrv12
    port map (
            O => \N__63799\,
            I => comm_state_2
        );

    \I__15928\ : CascadeMux
    port map (
            O => \N__63784\,
            I => \N__63774\
        );

    \I__15927\ : InMux
    port map (
            O => \N__63783\,
            I => \N__63771\
        );

    \I__15926\ : CascadeMux
    port map (
            O => \N__63782\,
            I => \N__63757\
        );

    \I__15925\ : CascadeMux
    port map (
            O => \N__63781\,
            I => \N__63753\
        );

    \I__15924\ : CascadeMux
    port map (
            O => \N__63780\,
            I => \N__63749\
        );

    \I__15923\ : CascadeMux
    port map (
            O => \N__63779\,
            I => \N__63745\
        );

    \I__15922\ : InMux
    port map (
            O => \N__63778\,
            I => \N__63732\
        );

    \I__15921\ : InMux
    port map (
            O => \N__63777\,
            I => \N__63727\
        );

    \I__15920\ : InMux
    port map (
            O => \N__63774\,
            I => \N__63727\
        );

    \I__15919\ : LocalMux
    port map (
            O => \N__63771\,
            I => \N__63719\
        );

    \I__15918\ : CascadeMux
    port map (
            O => \N__63770\,
            I => \N__63714\
        );

    \I__15917\ : CascadeMux
    port map (
            O => \N__63769\,
            I => \N__63711\
        );

    \I__15916\ : CascadeMux
    port map (
            O => \N__63768\,
            I => \N__63708\
        );

    \I__15915\ : CascadeMux
    port map (
            O => \N__63767\,
            I => \N__63705\
        );

    \I__15914\ : CascadeMux
    port map (
            O => \N__63766\,
            I => \N__63702\
        );

    \I__15913\ : CascadeMux
    port map (
            O => \N__63765\,
            I => \N__63699\
        );

    \I__15912\ : CascadeMux
    port map (
            O => \N__63764\,
            I => \N__63696\
        );

    \I__15911\ : CascadeMux
    port map (
            O => \N__63763\,
            I => \N__63693\
        );

    \I__15910\ : CascadeMux
    port map (
            O => \N__63762\,
            I => \N__63690\
        );

    \I__15909\ : InMux
    port map (
            O => \N__63761\,
            I => \N__63687\
        );

    \I__15908\ : InMux
    port map (
            O => \N__63760\,
            I => \N__63670\
        );

    \I__15907\ : InMux
    port map (
            O => \N__63757\,
            I => \N__63670\
        );

    \I__15906\ : InMux
    port map (
            O => \N__63756\,
            I => \N__63670\
        );

    \I__15905\ : InMux
    port map (
            O => \N__63753\,
            I => \N__63670\
        );

    \I__15904\ : InMux
    port map (
            O => \N__63752\,
            I => \N__63670\
        );

    \I__15903\ : InMux
    port map (
            O => \N__63749\,
            I => \N__63670\
        );

    \I__15902\ : InMux
    port map (
            O => \N__63748\,
            I => \N__63670\
        );

    \I__15901\ : InMux
    port map (
            O => \N__63745\,
            I => \N__63670\
        );

    \I__15900\ : InMux
    port map (
            O => \N__63744\,
            I => \N__63667\
        );

    \I__15899\ : InMux
    port map (
            O => \N__63743\,
            I => \N__63656\
        );

    \I__15898\ : InMux
    port map (
            O => \N__63742\,
            I => \N__63656\
        );

    \I__15897\ : InMux
    port map (
            O => \N__63741\,
            I => \N__63656\
        );

    \I__15896\ : InMux
    port map (
            O => \N__63740\,
            I => \N__63656\
        );

    \I__15895\ : InMux
    port map (
            O => \N__63739\,
            I => \N__63656\
        );

    \I__15894\ : InMux
    port map (
            O => \N__63738\,
            I => \N__63651\
        );

    \I__15893\ : CascadeMux
    port map (
            O => \N__63737\,
            I => \N__63645\
        );

    \I__15892\ : InMux
    port map (
            O => \N__63736\,
            I => \N__63637\
        );

    \I__15891\ : InMux
    port map (
            O => \N__63735\,
            I => \N__63637\
        );

    \I__15890\ : LocalMux
    port map (
            O => \N__63732\,
            I => \N__63634\
        );

    \I__15889\ : LocalMux
    port map (
            O => \N__63727\,
            I => \N__63631\
        );

    \I__15888\ : InMux
    port map (
            O => \N__63726\,
            I => \N__63628\
        );

    \I__15887\ : InMux
    port map (
            O => \N__63725\,
            I => \N__63625\
        );

    \I__15886\ : InMux
    port map (
            O => \N__63724\,
            I => \N__63622\
        );

    \I__15885\ : CascadeMux
    port map (
            O => \N__63723\,
            I => \N__63619\
        );

    \I__15884\ : InMux
    port map (
            O => \N__63722\,
            I => \N__63614\
        );

    \I__15883\ : Span4Mux_v
    port map (
            O => \N__63719\,
            I => \N__63598\
        );

    \I__15882\ : InMux
    port map (
            O => \N__63718\,
            I => \N__63589\
        );

    \I__15881\ : InMux
    port map (
            O => \N__63717\,
            I => \N__63589\
        );

    \I__15880\ : InMux
    port map (
            O => \N__63714\,
            I => \N__63580\
        );

    \I__15879\ : InMux
    port map (
            O => \N__63711\,
            I => \N__63580\
        );

    \I__15878\ : InMux
    port map (
            O => \N__63708\,
            I => \N__63580\
        );

    \I__15877\ : InMux
    port map (
            O => \N__63705\,
            I => \N__63580\
        );

    \I__15876\ : InMux
    port map (
            O => \N__63702\,
            I => \N__63571\
        );

    \I__15875\ : InMux
    port map (
            O => \N__63699\,
            I => \N__63571\
        );

    \I__15874\ : InMux
    port map (
            O => \N__63696\,
            I => \N__63571\
        );

    \I__15873\ : InMux
    port map (
            O => \N__63693\,
            I => \N__63571\
        );

    \I__15872\ : InMux
    port map (
            O => \N__63690\,
            I => \N__63568\
        );

    \I__15871\ : LocalMux
    port map (
            O => \N__63687\,
            I => \N__63559\
        );

    \I__15870\ : LocalMux
    port map (
            O => \N__63670\,
            I => \N__63559\
        );

    \I__15869\ : LocalMux
    port map (
            O => \N__63667\,
            I => \N__63559\
        );

    \I__15868\ : LocalMux
    port map (
            O => \N__63656\,
            I => \N__63559\
        );

    \I__15867\ : InMux
    port map (
            O => \N__63655\,
            I => \N__63554\
        );

    \I__15866\ : InMux
    port map (
            O => \N__63654\,
            I => \N__63554\
        );

    \I__15865\ : LocalMux
    port map (
            O => \N__63651\,
            I => \N__63551\
        );

    \I__15864\ : InMux
    port map (
            O => \N__63650\,
            I => \N__63548\
        );

    \I__15863\ : InMux
    port map (
            O => \N__63649\,
            I => \N__63545\
        );

    \I__15862\ : InMux
    port map (
            O => \N__63648\,
            I => \N__63542\
        );

    \I__15861\ : InMux
    port map (
            O => \N__63645\,
            I => \N__63536\
        );

    \I__15860\ : InMux
    port map (
            O => \N__63644\,
            I => \N__63529\
        );

    \I__15859\ : InMux
    port map (
            O => \N__63643\,
            I => \N__63529\
        );

    \I__15858\ : InMux
    port map (
            O => \N__63642\,
            I => \N__63529\
        );

    \I__15857\ : LocalMux
    port map (
            O => \N__63637\,
            I => \N__63514\
        );

    \I__15856\ : Span4Mux_h
    port map (
            O => \N__63634\,
            I => \N__63514\
        );

    \I__15855\ : Span4Mux_v
    port map (
            O => \N__63631\,
            I => \N__63514\
        );

    \I__15854\ : LocalMux
    port map (
            O => \N__63628\,
            I => \N__63514\
        );

    \I__15853\ : LocalMux
    port map (
            O => \N__63625\,
            I => \N__63514\
        );

    \I__15852\ : LocalMux
    port map (
            O => \N__63622\,
            I => \N__63511\
        );

    \I__15851\ : InMux
    port map (
            O => \N__63619\,
            I => \N__63506\
        );

    \I__15850\ : InMux
    port map (
            O => \N__63618\,
            I => \N__63506\
        );

    \I__15849\ : SRMux
    port map (
            O => \N__63617\,
            I => \N__63501\
        );

    \I__15848\ : LocalMux
    port map (
            O => \N__63614\,
            I => \N__63498\
        );

    \I__15847\ : InMux
    port map (
            O => \N__63613\,
            I => \N__63495\
        );

    \I__15846\ : InMux
    port map (
            O => \N__63612\,
            I => \N__63479\
        );

    \I__15845\ : InMux
    port map (
            O => \N__63611\,
            I => \N__63474\
        );

    \I__15844\ : InMux
    port map (
            O => \N__63610\,
            I => \N__63474\
        );

    \I__15843\ : InMux
    port map (
            O => \N__63609\,
            I => \N__63469\
        );

    \I__15842\ : InMux
    port map (
            O => \N__63608\,
            I => \N__63469\
        );

    \I__15841\ : InMux
    port map (
            O => \N__63607\,
            I => \N__63466\
        );

    \I__15840\ : InMux
    port map (
            O => \N__63606\,
            I => \N__63457\
        );

    \I__15839\ : InMux
    port map (
            O => \N__63605\,
            I => \N__63457\
        );

    \I__15838\ : InMux
    port map (
            O => \N__63604\,
            I => \N__63457\
        );

    \I__15837\ : InMux
    port map (
            O => \N__63603\,
            I => \N__63457\
        );

    \I__15836\ : InMux
    port map (
            O => \N__63602\,
            I => \N__63454\
        );

    \I__15835\ : InMux
    port map (
            O => \N__63601\,
            I => \N__63451\
        );

    \I__15834\ : Span4Mux_h
    port map (
            O => \N__63598\,
            I => \N__63448\
        );

    \I__15833\ : InMux
    port map (
            O => \N__63597\,
            I => \N__63445\
        );

    \I__15832\ : InMux
    port map (
            O => \N__63596\,
            I => \N__63438\
        );

    \I__15831\ : InMux
    port map (
            O => \N__63595\,
            I => \N__63438\
        );

    \I__15830\ : InMux
    port map (
            O => \N__63594\,
            I => \N__63438\
        );

    \I__15829\ : LocalMux
    port map (
            O => \N__63589\,
            I => \N__63421\
        );

    \I__15828\ : LocalMux
    port map (
            O => \N__63580\,
            I => \N__63421\
        );

    \I__15827\ : LocalMux
    port map (
            O => \N__63571\,
            I => \N__63421\
        );

    \I__15826\ : LocalMux
    port map (
            O => \N__63568\,
            I => \N__63421\
        );

    \I__15825\ : Span4Mux_v
    port map (
            O => \N__63559\,
            I => \N__63421\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__63554\,
            I => \N__63421\
        );

    \I__15823\ : Span4Mux_v
    port map (
            O => \N__63551\,
            I => \N__63421\
        );

    \I__15822\ : LocalMux
    port map (
            O => \N__63548\,
            I => \N__63421\
        );

    \I__15821\ : LocalMux
    port map (
            O => \N__63545\,
            I => \N__63418\
        );

    \I__15820\ : LocalMux
    port map (
            O => \N__63542\,
            I => \N__63415\
        );

    \I__15819\ : InMux
    port map (
            O => \N__63541\,
            I => \N__63412\
        );

    \I__15818\ : InMux
    port map (
            O => \N__63540\,
            I => \N__63407\
        );

    \I__15817\ : InMux
    port map (
            O => \N__63539\,
            I => \N__63407\
        );

    \I__15816\ : LocalMux
    port map (
            O => \N__63536\,
            I => \N__63402\
        );

    \I__15815\ : LocalMux
    port map (
            O => \N__63529\,
            I => \N__63402\
        );

    \I__15814\ : InMux
    port map (
            O => \N__63528\,
            I => \N__63397\
        );

    \I__15813\ : InMux
    port map (
            O => \N__63527\,
            I => \N__63397\
        );

    \I__15812\ : InMux
    port map (
            O => \N__63526\,
            I => \N__63394\
        );

    \I__15811\ : InMux
    port map (
            O => \N__63525\,
            I => \N__63390\
        );

    \I__15810\ : Span4Mux_v
    port map (
            O => \N__63514\,
            I => \N__63383\
        );

    \I__15809\ : Span4Mux_v
    port map (
            O => \N__63511\,
            I => \N__63383\
        );

    \I__15808\ : LocalMux
    port map (
            O => \N__63506\,
            I => \N__63383\
        );

    \I__15807\ : InMux
    port map (
            O => \N__63505\,
            I => \N__63373\
        );

    \I__15806\ : InMux
    port map (
            O => \N__63504\,
            I => \N__63373\
        );

    \I__15805\ : LocalMux
    port map (
            O => \N__63501\,
            I => \N__63366\
        );

    \I__15804\ : Span4Mux_h
    port map (
            O => \N__63498\,
            I => \N__63366\
        );

    \I__15803\ : LocalMux
    port map (
            O => \N__63495\,
            I => \N__63366\
        );

    \I__15802\ : InMux
    port map (
            O => \N__63494\,
            I => \N__63359\
        );

    \I__15801\ : InMux
    port map (
            O => \N__63493\,
            I => \N__63359\
        );

    \I__15800\ : InMux
    port map (
            O => \N__63492\,
            I => \N__63359\
        );

    \I__15799\ : InMux
    port map (
            O => \N__63491\,
            I => \N__63354\
        );

    \I__15798\ : InMux
    port map (
            O => \N__63490\,
            I => \N__63349\
        );

    \I__15797\ : InMux
    port map (
            O => \N__63489\,
            I => \N__63349\
        );

    \I__15796\ : InMux
    port map (
            O => \N__63488\,
            I => \N__63346\
        );

    \I__15795\ : InMux
    port map (
            O => \N__63487\,
            I => \N__63341\
        );

    \I__15794\ : InMux
    port map (
            O => \N__63486\,
            I => \N__63341\
        );

    \I__15793\ : InMux
    port map (
            O => \N__63485\,
            I => \N__63338\
        );

    \I__15792\ : InMux
    port map (
            O => \N__63484\,
            I => \N__63331\
        );

    \I__15791\ : InMux
    port map (
            O => \N__63483\,
            I => \N__63331\
        );

    \I__15790\ : InMux
    port map (
            O => \N__63482\,
            I => \N__63331\
        );

    \I__15789\ : LocalMux
    port map (
            O => \N__63479\,
            I => \N__63320\
        );

    \I__15788\ : LocalMux
    port map (
            O => \N__63474\,
            I => \N__63320\
        );

    \I__15787\ : LocalMux
    port map (
            O => \N__63469\,
            I => \N__63320\
        );

    \I__15786\ : LocalMux
    port map (
            O => \N__63466\,
            I => \N__63320\
        );

    \I__15785\ : LocalMux
    port map (
            O => \N__63457\,
            I => \N__63320\
        );

    \I__15784\ : LocalMux
    port map (
            O => \N__63454\,
            I => \N__63317\
        );

    \I__15783\ : LocalMux
    port map (
            O => \N__63451\,
            I => \N__63314\
        );

    \I__15782\ : Span4Mux_h
    port map (
            O => \N__63448\,
            I => \N__63305\
        );

    \I__15781\ : LocalMux
    port map (
            O => \N__63445\,
            I => \N__63305\
        );

    \I__15780\ : LocalMux
    port map (
            O => \N__63438\,
            I => \N__63305\
        );

    \I__15779\ : Span4Mux_v
    port map (
            O => \N__63421\,
            I => \N__63305\
        );

    \I__15778\ : Span4Mux_v
    port map (
            O => \N__63418\,
            I => \N__63300\
        );

    \I__15777\ : Span4Mux_v
    port map (
            O => \N__63415\,
            I => \N__63300\
        );

    \I__15776\ : LocalMux
    port map (
            O => \N__63412\,
            I => \N__63291\
        );

    \I__15775\ : LocalMux
    port map (
            O => \N__63407\,
            I => \N__63291\
        );

    \I__15774\ : Span4Mux_v
    port map (
            O => \N__63402\,
            I => \N__63291\
        );

    \I__15773\ : LocalMux
    port map (
            O => \N__63397\,
            I => \N__63291\
        );

    \I__15772\ : LocalMux
    port map (
            O => \N__63394\,
            I => \N__63288\
        );

    \I__15771\ : InMux
    port map (
            O => \N__63393\,
            I => \N__63285\
        );

    \I__15770\ : LocalMux
    port map (
            O => \N__63390\,
            I => \N__63282\
        );

    \I__15769\ : Span4Mux_h
    port map (
            O => \N__63383\,
            I => \N__63279\
        );

    \I__15768\ : InMux
    port map (
            O => \N__63382\,
            I => \N__63270\
        );

    \I__15767\ : InMux
    port map (
            O => \N__63381\,
            I => \N__63270\
        );

    \I__15766\ : InMux
    port map (
            O => \N__63380\,
            I => \N__63270\
        );

    \I__15765\ : InMux
    port map (
            O => \N__63379\,
            I => \N__63270\
        );

    \I__15764\ : InMux
    port map (
            O => \N__63378\,
            I => \N__63267\
        );

    \I__15763\ : LocalMux
    port map (
            O => \N__63373\,
            I => \N__63260\
        );

    \I__15762\ : Span4Mux_h
    port map (
            O => \N__63366\,
            I => \N__63260\
        );

    \I__15761\ : LocalMux
    port map (
            O => \N__63359\,
            I => \N__63260\
        );

    \I__15760\ : InMux
    port map (
            O => \N__63358\,
            I => \N__63255\
        );

    \I__15759\ : InMux
    port map (
            O => \N__63357\,
            I => \N__63255\
        );

    \I__15758\ : LocalMux
    port map (
            O => \N__63354\,
            I => \N__63240\
        );

    \I__15757\ : LocalMux
    port map (
            O => \N__63349\,
            I => \N__63240\
        );

    \I__15756\ : LocalMux
    port map (
            O => \N__63346\,
            I => \N__63240\
        );

    \I__15755\ : LocalMux
    port map (
            O => \N__63341\,
            I => \N__63240\
        );

    \I__15754\ : LocalMux
    port map (
            O => \N__63338\,
            I => \N__63240\
        );

    \I__15753\ : LocalMux
    port map (
            O => \N__63331\,
            I => \N__63240\
        );

    \I__15752\ : Span12Mux_v
    port map (
            O => \N__63320\,
            I => \N__63240\
        );

    \I__15751\ : Span4Mux_v
    port map (
            O => \N__63317\,
            I => \N__63229\
        );

    \I__15750\ : Span4Mux_v
    port map (
            O => \N__63314\,
            I => \N__63229\
        );

    \I__15749\ : Span4Mux_v
    port map (
            O => \N__63305\,
            I => \N__63229\
        );

    \I__15748\ : Span4Mux_h
    port map (
            O => \N__63300\,
            I => \N__63229\
        );

    \I__15747\ : Span4Mux_v
    port map (
            O => \N__63291\,
            I => \N__63229\
        );

    \I__15746\ : Span12Mux_h
    port map (
            O => \N__63288\,
            I => \N__63218\
        );

    \I__15745\ : LocalMux
    port map (
            O => \N__63285\,
            I => \N__63218\
        );

    \I__15744\ : Span12Mux_s9_v
    port map (
            O => \N__63282\,
            I => \N__63218\
        );

    \I__15743\ : Sp12to4
    port map (
            O => \N__63279\,
            I => \N__63218\
        );

    \I__15742\ : LocalMux
    port map (
            O => \N__63270\,
            I => \N__63218\
        );

    \I__15741\ : LocalMux
    port map (
            O => \N__63267\,
            I => comm_state_3
        );

    \I__15740\ : Odrv4
    port map (
            O => \N__63260\,
            I => comm_state_3
        );

    \I__15739\ : LocalMux
    port map (
            O => \N__63255\,
            I => comm_state_3
        );

    \I__15738\ : Odrv12
    port map (
            O => \N__63240\,
            I => comm_state_3
        );

    \I__15737\ : Odrv4
    port map (
            O => \N__63229\,
            I => comm_state_3
        );

    \I__15736\ : Odrv12
    port map (
            O => \N__63218\,
            I => comm_state_3
        );

    \I__15735\ : CascadeMux
    port map (
            O => \N__63205\,
            I => \N__63201\
        );

    \I__15734\ : InMux
    port map (
            O => \N__63204\,
            I => \N__63197\
        );

    \I__15733\ : InMux
    port map (
            O => \N__63201\,
            I => \N__63191\
        );

    \I__15732\ : CascadeMux
    port map (
            O => \N__63200\,
            I => \N__63185\
        );

    \I__15731\ : LocalMux
    port map (
            O => \N__63197\,
            I => \N__63182\
        );

    \I__15730\ : InMux
    port map (
            O => \N__63196\,
            I => \N__63177\
        );

    \I__15729\ : InMux
    port map (
            O => \N__63195\,
            I => \N__63177\
        );

    \I__15728\ : InMux
    port map (
            O => \N__63194\,
            I => \N__63174\
        );

    \I__15727\ : LocalMux
    port map (
            O => \N__63191\,
            I => \N__63170\
        );

    \I__15726\ : InMux
    port map (
            O => \N__63190\,
            I => \N__63167\
        );

    \I__15725\ : CascadeMux
    port map (
            O => \N__63189\,
            I => \N__63164\
        );

    \I__15724\ : InMux
    port map (
            O => \N__63188\,
            I => \N__63157\
        );

    \I__15723\ : InMux
    port map (
            O => \N__63185\,
            I => \N__63157\
        );

    \I__15722\ : Span4Mux_v
    port map (
            O => \N__63182\,
            I => \N__63152\
        );

    \I__15721\ : LocalMux
    port map (
            O => \N__63177\,
            I => \N__63152\
        );

    \I__15720\ : LocalMux
    port map (
            O => \N__63174\,
            I => \N__63149\
        );

    \I__15719\ : InMux
    port map (
            O => \N__63173\,
            I => \N__63146\
        );

    \I__15718\ : Span4Mux_v
    port map (
            O => \N__63170\,
            I => \N__63140\
        );

    \I__15717\ : LocalMux
    port map (
            O => \N__63167\,
            I => \N__63140\
        );

    \I__15716\ : InMux
    port map (
            O => \N__63164\,
            I => \N__63133\
        );

    \I__15715\ : InMux
    port map (
            O => \N__63163\,
            I => \N__63133\
        );

    \I__15714\ : InMux
    port map (
            O => \N__63162\,
            I => \N__63133\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__63157\,
            I => \N__63128\
        );

    \I__15712\ : Span4Mux_v
    port map (
            O => \N__63152\,
            I => \N__63128\
        );

    \I__15711\ : Span4Mux_h
    port map (
            O => \N__63149\,
            I => \N__63125\
        );

    \I__15710\ : LocalMux
    port map (
            O => \N__63146\,
            I => \N__63122\
        );

    \I__15709\ : InMux
    port map (
            O => \N__63145\,
            I => \N__63119\
        );

    \I__15708\ : Span4Mux_h
    port map (
            O => \N__63140\,
            I => \N__63114\
        );

    \I__15707\ : LocalMux
    port map (
            O => \N__63133\,
            I => \N__63114\
        );

    \I__15706\ : Span4Mux_v
    port map (
            O => \N__63128\,
            I => \N__63111\
        );

    \I__15705\ : Span4Mux_v
    port map (
            O => \N__63125\,
            I => \N__63105\
        );

    \I__15704\ : Span4Mux_v
    port map (
            O => \N__63122\,
            I => \N__63105\
        );

    \I__15703\ : LocalMux
    port map (
            O => \N__63119\,
            I => \N__63100\
        );

    \I__15702\ : Span4Mux_h
    port map (
            O => \N__63114\,
            I => \N__63100\
        );

    \I__15701\ : Sp12to4
    port map (
            O => \N__63111\,
            I => \N__63097\
        );

    \I__15700\ : InMux
    port map (
            O => \N__63110\,
            I => \N__63094\
        );

    \I__15699\ : Odrv4
    port map (
            O => \N__63105\,
            I => n12966
        );

    \I__15698\ : Odrv4
    port map (
            O => \N__63100\,
            I => n12966
        );

    \I__15697\ : Odrv12
    port map (
            O => \N__63097\,
            I => n12966
        );

    \I__15696\ : LocalMux
    port map (
            O => \N__63094\,
            I => n12966
        );

    \I__15695\ : CascadeMux
    port map (
            O => \N__63085\,
            I => \N__63067\
        );

    \I__15694\ : InMux
    port map (
            O => \N__63084\,
            I => \N__63061\
        );

    \I__15693\ : InMux
    port map (
            O => \N__63083\,
            I => \N__63061\
        );

    \I__15692\ : InMux
    port map (
            O => \N__63082\,
            I => \N__63052\
        );

    \I__15691\ : InMux
    port map (
            O => \N__63081\,
            I => \N__63042\
        );

    \I__15690\ : InMux
    port map (
            O => \N__63080\,
            I => \N__63039\
        );

    \I__15689\ : InMux
    port map (
            O => \N__63079\,
            I => \N__63034\
        );

    \I__15688\ : InMux
    port map (
            O => \N__63078\,
            I => \N__63034\
        );

    \I__15687\ : InMux
    port map (
            O => \N__63077\,
            I => \N__63031\
        );

    \I__15686\ : InMux
    port map (
            O => \N__63076\,
            I => \N__63024\
        );

    \I__15685\ : CascadeMux
    port map (
            O => \N__63075\,
            I => \N__63021\
        );

    \I__15684\ : InMux
    port map (
            O => \N__63074\,
            I => \N__63018\
        );

    \I__15683\ : InMux
    port map (
            O => \N__63073\,
            I => \N__63015\
        );

    \I__15682\ : InMux
    port map (
            O => \N__63072\,
            I => \N__63012\
        );

    \I__15681\ : InMux
    port map (
            O => \N__63071\,
            I => \N__63003\
        );

    \I__15680\ : InMux
    port map (
            O => \N__63070\,
            I => \N__63003\
        );

    \I__15679\ : InMux
    port map (
            O => \N__63067\,
            I => \N__63003\
        );

    \I__15678\ : InMux
    port map (
            O => \N__63066\,
            I => \N__63003\
        );

    \I__15677\ : LocalMux
    port map (
            O => \N__63061\,
            I => \N__63000\
        );

    \I__15676\ : InMux
    port map (
            O => \N__63060\,
            I => \N__62991\
        );

    \I__15675\ : InMux
    port map (
            O => \N__63059\,
            I => \N__62991\
        );

    \I__15674\ : InMux
    port map (
            O => \N__63058\,
            I => \N__62991\
        );

    \I__15673\ : InMux
    port map (
            O => \N__63057\,
            I => \N__62991\
        );

    \I__15672\ : InMux
    port map (
            O => \N__63056\,
            I => \N__62986\
        );

    \I__15671\ : InMux
    port map (
            O => \N__63055\,
            I => \N__62986\
        );

    \I__15670\ : LocalMux
    port map (
            O => \N__63052\,
            I => \N__62983\
        );

    \I__15669\ : InMux
    port map (
            O => \N__63051\,
            I => \N__62980\
        );

    \I__15668\ : InMux
    port map (
            O => \N__63050\,
            I => \N__62973\
        );

    \I__15667\ : InMux
    port map (
            O => \N__63049\,
            I => \N__62973\
        );

    \I__15666\ : InMux
    port map (
            O => \N__63048\,
            I => \N__62973\
        );

    \I__15665\ : InMux
    port map (
            O => \N__63047\,
            I => \N__62970\
        );

    \I__15664\ : InMux
    port map (
            O => \N__63046\,
            I => \N__62964\
        );

    \I__15663\ : InMux
    port map (
            O => \N__63045\,
            I => \N__62964\
        );

    \I__15662\ : LocalMux
    port map (
            O => \N__63042\,
            I => \N__62957\
        );

    \I__15661\ : LocalMux
    port map (
            O => \N__63039\,
            I => \N__62957\
        );

    \I__15660\ : LocalMux
    port map (
            O => \N__63034\,
            I => \N__62957\
        );

    \I__15659\ : LocalMux
    port map (
            O => \N__63031\,
            I => \N__62954\
        );

    \I__15658\ : InMux
    port map (
            O => \N__63030\,
            I => \N__62949\
        );

    \I__15657\ : InMux
    port map (
            O => \N__63029\,
            I => \N__62949\
        );

    \I__15656\ : InMux
    port map (
            O => \N__63028\,
            I => \N__62944\
        );

    \I__15655\ : InMux
    port map (
            O => \N__63027\,
            I => \N__62944\
        );

    \I__15654\ : LocalMux
    port map (
            O => \N__63024\,
            I => \N__62940\
        );

    \I__15653\ : InMux
    port map (
            O => \N__63021\,
            I => \N__62937\
        );

    \I__15652\ : LocalMux
    port map (
            O => \N__63018\,
            I => \N__62927\
        );

    \I__15651\ : LocalMux
    port map (
            O => \N__63015\,
            I => \N__62924\
        );

    \I__15650\ : LocalMux
    port map (
            O => \N__63012\,
            I => \N__62913\
        );

    \I__15649\ : LocalMux
    port map (
            O => \N__63003\,
            I => \N__62913\
        );

    \I__15648\ : Span4Mux_v
    port map (
            O => \N__63000\,
            I => \N__62913\
        );

    \I__15647\ : LocalMux
    port map (
            O => \N__62991\,
            I => \N__62913\
        );

    \I__15646\ : LocalMux
    port map (
            O => \N__62986\,
            I => \N__62913\
        );

    \I__15645\ : Span4Mux_v
    port map (
            O => \N__62983\,
            I => \N__62908\
        );

    \I__15644\ : LocalMux
    port map (
            O => \N__62980\,
            I => \N__62908\
        );

    \I__15643\ : LocalMux
    port map (
            O => \N__62973\,
            I => \N__62902\
        );

    \I__15642\ : LocalMux
    port map (
            O => \N__62970\,
            I => \N__62899\
        );

    \I__15641\ : InMux
    port map (
            O => \N__62969\,
            I => \N__62896\
        );

    \I__15640\ : LocalMux
    port map (
            O => \N__62964\,
            I => \N__62891\
        );

    \I__15639\ : Span4Mux_v
    port map (
            O => \N__62957\,
            I => \N__62891\
        );

    \I__15638\ : Span4Mux_h
    port map (
            O => \N__62954\,
            I => \N__62884\
        );

    \I__15637\ : LocalMux
    port map (
            O => \N__62949\,
            I => \N__62884\
        );

    \I__15636\ : LocalMux
    port map (
            O => \N__62944\,
            I => \N__62884\
        );

    \I__15635\ : InMux
    port map (
            O => \N__62943\,
            I => \N__62881\
        );

    \I__15634\ : Span4Mux_h
    port map (
            O => \N__62940\,
            I => \N__62878\
        );

    \I__15633\ : LocalMux
    port map (
            O => \N__62937\,
            I => \N__62875\
        );

    \I__15632\ : InMux
    port map (
            O => \N__62936\,
            I => \N__62872\
        );

    \I__15631\ : InMux
    port map (
            O => \N__62935\,
            I => \N__62863\
        );

    \I__15630\ : InMux
    port map (
            O => \N__62934\,
            I => \N__62863\
        );

    \I__15629\ : InMux
    port map (
            O => \N__62933\,
            I => \N__62863\
        );

    \I__15628\ : InMux
    port map (
            O => \N__62932\,
            I => \N__62863\
        );

    \I__15627\ : InMux
    port map (
            O => \N__62931\,
            I => \N__62858\
        );

    \I__15626\ : InMux
    port map (
            O => \N__62930\,
            I => \N__62858\
        );

    \I__15625\ : Span4Mux_h
    port map (
            O => \N__62927\,
            I => \N__62849\
        );

    \I__15624\ : Span4Mux_v
    port map (
            O => \N__62924\,
            I => \N__62849\
        );

    \I__15623\ : Span4Mux_v
    port map (
            O => \N__62913\,
            I => \N__62849\
        );

    \I__15622\ : Span4Mux_v
    port map (
            O => \N__62908\,
            I => \N__62849\
        );

    \I__15621\ : InMux
    port map (
            O => \N__62907\,
            I => \N__62844\
        );

    \I__15620\ : InMux
    port map (
            O => \N__62906\,
            I => \N__62844\
        );

    \I__15619\ : InMux
    port map (
            O => \N__62905\,
            I => \N__62841\
        );

    \I__15618\ : Sp12to4
    port map (
            O => \N__62902\,
            I => \N__62836\
        );

    \I__15617\ : Span12Mux_h
    port map (
            O => \N__62899\,
            I => \N__62836\
        );

    \I__15616\ : LocalMux
    port map (
            O => \N__62896\,
            I => \N__62831\
        );

    \I__15615\ : Span4Mux_h
    port map (
            O => \N__62891\,
            I => \N__62831\
        );

    \I__15614\ : Span4Mux_h
    port map (
            O => \N__62884\,
            I => \N__62822\
        );

    \I__15613\ : LocalMux
    port map (
            O => \N__62881\,
            I => \N__62822\
        );

    \I__15612\ : Span4Mux_h
    port map (
            O => \N__62878\,
            I => \N__62822\
        );

    \I__15611\ : Span4Mux_h
    port map (
            O => \N__62875\,
            I => \N__62822\
        );

    \I__15610\ : LocalMux
    port map (
            O => \N__62872\,
            I => comm_state_0
        );

    \I__15609\ : LocalMux
    port map (
            O => \N__62863\,
            I => comm_state_0
        );

    \I__15608\ : LocalMux
    port map (
            O => \N__62858\,
            I => comm_state_0
        );

    \I__15607\ : Odrv4
    port map (
            O => \N__62849\,
            I => comm_state_0
        );

    \I__15606\ : LocalMux
    port map (
            O => \N__62844\,
            I => comm_state_0
        );

    \I__15605\ : LocalMux
    port map (
            O => \N__62841\,
            I => comm_state_0
        );

    \I__15604\ : Odrv12
    port map (
            O => \N__62836\,
            I => comm_state_0
        );

    \I__15603\ : Odrv4
    port map (
            O => \N__62831\,
            I => comm_state_0
        );

    \I__15602\ : Odrv4
    port map (
            O => \N__62822\,
            I => comm_state_0
        );

    \I__15601\ : CEMux
    port map (
            O => \N__62803\,
            I => \N__62800\
        );

    \I__15600\ : LocalMux
    port map (
            O => \N__62800\,
            I => \N__62797\
        );

    \I__15599\ : Odrv4
    port map (
            O => \N__62797\,
            I => n12045
        );

    \I__15598\ : CascadeMux
    port map (
            O => \N__62794\,
            I => \N__62791\
        );

    \I__15597\ : InMux
    port map (
            O => \N__62791\,
            I => \N__62785\
        );

    \I__15596\ : InMux
    port map (
            O => \N__62790\,
            I => \N__62781\
        );

    \I__15595\ : InMux
    port map (
            O => \N__62789\,
            I => \N__62776\
        );

    \I__15594\ : InMux
    port map (
            O => \N__62788\,
            I => \N__62772\
        );

    \I__15593\ : LocalMux
    port map (
            O => \N__62785\,
            I => \N__62769\
        );

    \I__15592\ : InMux
    port map (
            O => \N__62784\,
            I => \N__62766\
        );

    \I__15591\ : LocalMux
    port map (
            O => \N__62781\,
            I => \N__62763\
        );

    \I__15590\ : InMux
    port map (
            O => \N__62780\,
            I => \N__62760\
        );

    \I__15589\ : CascadeMux
    port map (
            O => \N__62779\,
            I => \N__62757\
        );

    \I__15588\ : LocalMux
    port map (
            O => \N__62776\,
            I => \N__62754\
        );

    \I__15587\ : CascadeMux
    port map (
            O => \N__62775\,
            I => \N__62751\
        );

    \I__15586\ : LocalMux
    port map (
            O => \N__62772\,
            I => \N__62748\
        );

    \I__15585\ : Span4Mux_v
    port map (
            O => \N__62769\,
            I => \N__62743\
        );

    \I__15584\ : LocalMux
    port map (
            O => \N__62766\,
            I => \N__62743\
        );

    \I__15583\ : Span4Mux_v
    port map (
            O => \N__62763\,
            I => \N__62740\
        );

    \I__15582\ : LocalMux
    port map (
            O => \N__62760\,
            I => \N__62737\
        );

    \I__15581\ : InMux
    port map (
            O => \N__62757\,
            I => \N__62734\
        );

    \I__15580\ : Span4Mux_h
    port map (
            O => \N__62754\,
            I => \N__62731\
        );

    \I__15579\ : InMux
    port map (
            O => \N__62751\,
            I => \N__62728\
        );

    \I__15578\ : Span4Mux_h
    port map (
            O => \N__62748\,
            I => \N__62724\
        );

    \I__15577\ : Span4Mux_v
    port map (
            O => \N__62743\,
            I => \N__62721\
        );

    \I__15576\ : Span4Mux_h
    port map (
            O => \N__62740\,
            I => \N__62716\
        );

    \I__15575\ : Span4Mux_v
    port map (
            O => \N__62737\,
            I => \N__62716\
        );

    \I__15574\ : LocalMux
    port map (
            O => \N__62734\,
            I => \N__62713\
        );

    \I__15573\ : Span4Mux_h
    port map (
            O => \N__62731\,
            I => \N__62708\
        );

    \I__15572\ : LocalMux
    port map (
            O => \N__62728\,
            I => \N__62708\
        );

    \I__15571\ : InMux
    port map (
            O => \N__62727\,
            I => \N__62705\
        );

    \I__15570\ : Odrv4
    port map (
            O => \N__62724\,
            I => comm_rx_buf_3
        );

    \I__15569\ : Odrv4
    port map (
            O => \N__62721\,
            I => comm_rx_buf_3
        );

    \I__15568\ : Odrv4
    port map (
            O => \N__62716\,
            I => comm_rx_buf_3
        );

    \I__15567\ : Odrv12
    port map (
            O => \N__62713\,
            I => comm_rx_buf_3
        );

    \I__15566\ : Odrv4
    port map (
            O => \N__62708\,
            I => comm_rx_buf_3
        );

    \I__15565\ : LocalMux
    port map (
            O => \N__62705\,
            I => comm_rx_buf_3
        );

    \I__15564\ : InMux
    port map (
            O => \N__62692\,
            I => \N__62686\
        );

    \I__15563\ : CascadeMux
    port map (
            O => \N__62691\,
            I => \N__62682\
        );

    \I__15562\ : CascadeMux
    port map (
            O => \N__62690\,
            I => \N__62679\
        );

    \I__15561\ : InMux
    port map (
            O => \N__62689\,
            I => \N__62667\
        );

    \I__15560\ : LocalMux
    port map (
            O => \N__62686\,
            I => \N__62664\
        );

    \I__15559\ : CascadeMux
    port map (
            O => \N__62685\,
            I => \N__62649\
        );

    \I__15558\ : InMux
    port map (
            O => \N__62682\,
            I => \N__62638\
        );

    \I__15557\ : InMux
    port map (
            O => \N__62679\,
            I => \N__62638\
        );

    \I__15556\ : InMux
    port map (
            O => \N__62678\,
            I => \N__62638\
        );

    \I__15555\ : CascadeMux
    port map (
            O => \N__62677\,
            I => \N__62634\
        );

    \I__15554\ : CascadeMux
    port map (
            O => \N__62676\,
            I => \N__62612\
        );

    \I__15553\ : InMux
    port map (
            O => \N__62675\,
            I => \N__62588\
        );

    \I__15552\ : InMux
    port map (
            O => \N__62674\,
            I => \N__62588\
        );

    \I__15551\ : InMux
    port map (
            O => \N__62673\,
            I => \N__62588\
        );

    \I__15550\ : InMux
    port map (
            O => \N__62672\,
            I => \N__62585\
        );

    \I__15549\ : InMux
    port map (
            O => \N__62671\,
            I => \N__62582\
        );

    \I__15548\ : InMux
    port map (
            O => \N__62670\,
            I => \N__62579\
        );

    \I__15547\ : LocalMux
    port map (
            O => \N__62667\,
            I => \N__62576\
        );

    \I__15546\ : Span4Mux_v
    port map (
            O => \N__62664\,
            I => \N__62573\
        );

    \I__15545\ : InMux
    port map (
            O => \N__62663\,
            I => \N__62561\
        );

    \I__15544\ : InMux
    port map (
            O => \N__62662\,
            I => \N__62548\
        );

    \I__15543\ : InMux
    port map (
            O => \N__62661\,
            I => \N__62548\
        );

    \I__15542\ : InMux
    port map (
            O => \N__62660\,
            I => \N__62548\
        );

    \I__15541\ : InMux
    port map (
            O => \N__62659\,
            I => \N__62548\
        );

    \I__15540\ : InMux
    port map (
            O => \N__62658\,
            I => \N__62548\
        );

    \I__15539\ : InMux
    port map (
            O => \N__62657\,
            I => \N__62548\
        );

    \I__15538\ : InMux
    port map (
            O => \N__62656\,
            I => \N__62531\
        );

    \I__15537\ : InMux
    port map (
            O => \N__62655\,
            I => \N__62531\
        );

    \I__15536\ : InMux
    port map (
            O => \N__62654\,
            I => \N__62531\
        );

    \I__15535\ : InMux
    port map (
            O => \N__62653\,
            I => \N__62531\
        );

    \I__15534\ : InMux
    port map (
            O => \N__62652\,
            I => \N__62531\
        );

    \I__15533\ : InMux
    port map (
            O => \N__62649\,
            I => \N__62531\
        );

    \I__15532\ : InMux
    port map (
            O => \N__62648\,
            I => \N__62531\
        );

    \I__15531\ : InMux
    port map (
            O => \N__62647\,
            I => \N__62531\
        );

    \I__15530\ : InMux
    port map (
            O => \N__62646\,
            I => \N__62516\
        );

    \I__15529\ : InMux
    port map (
            O => \N__62645\,
            I => \N__62516\
        );

    \I__15528\ : LocalMux
    port map (
            O => \N__62638\,
            I => \N__62513\
        );

    \I__15527\ : InMux
    port map (
            O => \N__62637\,
            I => \N__62510\
        );

    \I__15526\ : InMux
    port map (
            O => \N__62634\,
            I => \N__62507\
        );

    \I__15525\ : CascadeMux
    port map (
            O => \N__62633\,
            I => \N__62504\
        );

    \I__15524\ : InMux
    port map (
            O => \N__62632\,
            I => \N__62487\
        );

    \I__15523\ : InMux
    port map (
            O => \N__62631\,
            I => \N__62487\
        );

    \I__15522\ : InMux
    port map (
            O => \N__62630\,
            I => \N__62487\
        );

    \I__15521\ : InMux
    port map (
            O => \N__62629\,
            I => \N__62487\
        );

    \I__15520\ : InMux
    port map (
            O => \N__62628\,
            I => \N__62487\
        );

    \I__15519\ : InMux
    port map (
            O => \N__62627\,
            I => \N__62487\
        );

    \I__15518\ : InMux
    port map (
            O => \N__62626\,
            I => \N__62487\
        );

    \I__15517\ : InMux
    port map (
            O => \N__62625\,
            I => \N__62487\
        );

    \I__15516\ : InMux
    port map (
            O => \N__62624\,
            I => \N__62482\
        );

    \I__15515\ : InMux
    port map (
            O => \N__62623\,
            I => \N__62463\
        );

    \I__15514\ : InMux
    port map (
            O => \N__62622\,
            I => \N__62463\
        );

    \I__15513\ : InMux
    port map (
            O => \N__62621\,
            I => \N__62463\
        );

    \I__15512\ : InMux
    port map (
            O => \N__62620\,
            I => \N__62463\
        );

    \I__15511\ : InMux
    port map (
            O => \N__62619\,
            I => \N__62463\
        );

    \I__15510\ : InMux
    port map (
            O => \N__62618\,
            I => \N__62463\
        );

    \I__15509\ : InMux
    port map (
            O => \N__62617\,
            I => \N__62463\
        );

    \I__15508\ : InMux
    port map (
            O => \N__62616\,
            I => \N__62463\
        );

    \I__15507\ : InMux
    port map (
            O => \N__62615\,
            I => \N__62460\
        );

    \I__15506\ : InMux
    port map (
            O => \N__62612\,
            I => \N__62451\
        );

    \I__15505\ : InMux
    port map (
            O => \N__62611\,
            I => \N__62451\
        );

    \I__15504\ : InMux
    port map (
            O => \N__62610\,
            I => \N__62451\
        );

    \I__15503\ : InMux
    port map (
            O => \N__62609\,
            I => \N__62451\
        );

    \I__15502\ : CascadeMux
    port map (
            O => \N__62608\,
            I => \N__62446\
        );

    \I__15501\ : InMux
    port map (
            O => \N__62607\,
            I => \N__62443\
        );

    \I__15500\ : InMux
    port map (
            O => \N__62606\,
            I => \N__62440\
        );

    \I__15499\ : InMux
    port map (
            O => \N__62605\,
            I => \N__62435\
        );

    \I__15498\ : InMux
    port map (
            O => \N__62604\,
            I => \N__62435\
        );

    \I__15497\ : InMux
    port map (
            O => \N__62603\,
            I => \N__62432\
        );

    \I__15496\ : InMux
    port map (
            O => \N__62602\,
            I => \N__62429\
        );

    \I__15495\ : CascadeMux
    port map (
            O => \N__62601\,
            I => \N__62423\
        );

    \I__15494\ : InMux
    port map (
            O => \N__62600\,
            I => \N__62418\
        );

    \I__15493\ : InMux
    port map (
            O => \N__62599\,
            I => \N__62411\
        );

    \I__15492\ : InMux
    port map (
            O => \N__62598\,
            I => \N__62411\
        );

    \I__15491\ : InMux
    port map (
            O => \N__62597\,
            I => \N__62411\
        );

    \I__15490\ : InMux
    port map (
            O => \N__62596\,
            I => \N__62406\
        );

    \I__15489\ : InMux
    port map (
            O => \N__62595\,
            I => \N__62406\
        );

    \I__15488\ : LocalMux
    port map (
            O => \N__62588\,
            I => \N__62403\
        );

    \I__15487\ : LocalMux
    port map (
            O => \N__62585\,
            I => \N__62392\
        );

    \I__15486\ : LocalMux
    port map (
            O => \N__62582\,
            I => \N__62392\
        );

    \I__15485\ : LocalMux
    port map (
            O => \N__62579\,
            I => \N__62392\
        );

    \I__15484\ : Span4Mux_h
    port map (
            O => \N__62576\,
            I => \N__62392\
        );

    \I__15483\ : Span4Mux_h
    port map (
            O => \N__62573\,
            I => \N__62392\
        );

    \I__15482\ : InMux
    port map (
            O => \N__62572\,
            I => \N__62385\
        );

    \I__15481\ : InMux
    port map (
            O => \N__62571\,
            I => \N__62385\
        );

    \I__15480\ : InMux
    port map (
            O => \N__62570\,
            I => \N__62385\
        );

    \I__15479\ : InMux
    port map (
            O => \N__62569\,
            I => \N__62380\
        );

    \I__15478\ : InMux
    port map (
            O => \N__62568\,
            I => \N__62380\
        );

    \I__15477\ : InMux
    port map (
            O => \N__62567\,
            I => \N__62373\
        );

    \I__15476\ : InMux
    port map (
            O => \N__62566\,
            I => \N__62373\
        );

    \I__15475\ : InMux
    port map (
            O => \N__62565\,
            I => \N__62373\
        );

    \I__15474\ : InMux
    port map (
            O => \N__62564\,
            I => \N__62370\
        );

    \I__15473\ : LocalMux
    port map (
            O => \N__62561\,
            I => \N__62361\
        );

    \I__15472\ : LocalMux
    port map (
            O => \N__62548\,
            I => \N__62361\
        );

    \I__15471\ : LocalMux
    port map (
            O => \N__62531\,
            I => \N__62361\
        );

    \I__15470\ : InMux
    port map (
            O => \N__62530\,
            I => \N__62358\
        );

    \I__15469\ : InMux
    port map (
            O => \N__62529\,
            I => \N__62355\
        );

    \I__15468\ : InMux
    port map (
            O => \N__62528\,
            I => \N__62338\
        );

    \I__15467\ : InMux
    port map (
            O => \N__62527\,
            I => \N__62338\
        );

    \I__15466\ : InMux
    port map (
            O => \N__62526\,
            I => \N__62338\
        );

    \I__15465\ : InMux
    port map (
            O => \N__62525\,
            I => \N__62338\
        );

    \I__15464\ : InMux
    port map (
            O => \N__62524\,
            I => \N__62338\
        );

    \I__15463\ : InMux
    port map (
            O => \N__62523\,
            I => \N__62338\
        );

    \I__15462\ : InMux
    port map (
            O => \N__62522\,
            I => \N__62338\
        );

    \I__15461\ : InMux
    port map (
            O => \N__62521\,
            I => \N__62338\
        );

    \I__15460\ : LocalMux
    port map (
            O => \N__62516\,
            I => \N__62335\
        );

    \I__15459\ : Span4Mux_v
    port map (
            O => \N__62513\,
            I => \N__62332\
        );

    \I__15458\ : LocalMux
    port map (
            O => \N__62510\,
            I => \N__62327\
        );

    \I__15457\ : LocalMux
    port map (
            O => \N__62507\,
            I => \N__62327\
        );

    \I__15456\ : InMux
    port map (
            O => \N__62504\,
            I => \N__62324\
        );

    \I__15455\ : LocalMux
    port map (
            O => \N__62487\,
            I => \N__62321\
        );

    \I__15454\ : InMux
    port map (
            O => \N__62486\,
            I => \N__62316\
        );

    \I__15453\ : InMux
    port map (
            O => \N__62485\,
            I => \N__62316\
        );

    \I__15452\ : LocalMux
    port map (
            O => \N__62482\,
            I => \N__62313\
        );

    \I__15451\ : InMux
    port map (
            O => \N__62481\,
            I => \N__62308\
        );

    \I__15450\ : InMux
    port map (
            O => \N__62480\,
            I => \N__62308\
        );

    \I__15449\ : LocalMux
    port map (
            O => \N__62463\,
            I => \N__62301\
        );

    \I__15448\ : LocalMux
    port map (
            O => \N__62460\,
            I => \N__62301\
        );

    \I__15447\ : LocalMux
    port map (
            O => \N__62451\,
            I => \N__62301\
        );

    \I__15446\ : InMux
    port map (
            O => \N__62450\,
            I => \N__62298\
        );

    \I__15445\ : InMux
    port map (
            O => \N__62449\,
            I => \N__62285\
        );

    \I__15444\ : InMux
    port map (
            O => \N__62446\,
            I => \N__62285\
        );

    \I__15443\ : LocalMux
    port map (
            O => \N__62443\,
            I => \N__62276\
        );

    \I__15442\ : LocalMux
    port map (
            O => \N__62440\,
            I => \N__62276\
        );

    \I__15441\ : LocalMux
    port map (
            O => \N__62435\,
            I => \N__62276\
        );

    \I__15440\ : LocalMux
    port map (
            O => \N__62432\,
            I => \N__62276\
        );

    \I__15439\ : LocalMux
    port map (
            O => \N__62429\,
            I => \N__62273\
        );

    \I__15438\ : InMux
    port map (
            O => \N__62428\,
            I => \N__62260\
        );

    \I__15437\ : InMux
    port map (
            O => \N__62427\,
            I => \N__62260\
        );

    \I__15436\ : InMux
    port map (
            O => \N__62426\,
            I => \N__62260\
        );

    \I__15435\ : InMux
    port map (
            O => \N__62423\,
            I => \N__62260\
        );

    \I__15434\ : InMux
    port map (
            O => \N__62422\,
            I => \N__62260\
        );

    \I__15433\ : InMux
    port map (
            O => \N__62421\,
            I => \N__62260\
        );

    \I__15432\ : LocalMux
    port map (
            O => \N__62418\,
            I => \N__62243\
        );

    \I__15431\ : LocalMux
    port map (
            O => \N__62411\,
            I => \N__62243\
        );

    \I__15430\ : LocalMux
    port map (
            O => \N__62406\,
            I => \N__62243\
        );

    \I__15429\ : Span4Mux_h
    port map (
            O => \N__62403\,
            I => \N__62243\
        );

    \I__15428\ : Span4Mux_v
    port map (
            O => \N__62392\,
            I => \N__62243\
        );

    \I__15427\ : LocalMux
    port map (
            O => \N__62385\,
            I => \N__62243\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__62380\,
            I => \N__62243\
        );

    \I__15425\ : LocalMux
    port map (
            O => \N__62373\,
            I => \N__62243\
        );

    \I__15424\ : LocalMux
    port map (
            O => \N__62370\,
            I => \N__62237\
        );

    \I__15423\ : InMux
    port map (
            O => \N__62369\,
            I => \N__62232\
        );

    \I__15422\ : InMux
    port map (
            O => \N__62368\,
            I => \N__62232\
        );

    \I__15421\ : Span4Mux_h
    port map (
            O => \N__62361\,
            I => \N__62227\
        );

    \I__15420\ : LocalMux
    port map (
            O => \N__62358\,
            I => \N__62227\
        );

    \I__15419\ : LocalMux
    port map (
            O => \N__62355\,
            I => \N__62218\
        );

    \I__15418\ : LocalMux
    port map (
            O => \N__62338\,
            I => \N__62218\
        );

    \I__15417\ : Span4Mux_v
    port map (
            O => \N__62335\,
            I => \N__62218\
        );

    \I__15416\ : Span4Mux_h
    port map (
            O => \N__62332\,
            I => \N__62218\
        );

    \I__15415\ : Span4Mux_h
    port map (
            O => \N__62327\,
            I => \N__62215\
        );

    \I__15414\ : LocalMux
    port map (
            O => \N__62324\,
            I => \N__62212\
        );

    \I__15413\ : Span4Mux_v
    port map (
            O => \N__62321\,
            I => \N__62205\
        );

    \I__15412\ : LocalMux
    port map (
            O => \N__62316\,
            I => \N__62205\
        );

    \I__15411\ : Span4Mux_h
    port map (
            O => \N__62313\,
            I => \N__62205\
        );

    \I__15410\ : LocalMux
    port map (
            O => \N__62308\,
            I => \N__62200\
        );

    \I__15409\ : Span4Mux_h
    port map (
            O => \N__62301\,
            I => \N__62200\
        );

    \I__15408\ : LocalMux
    port map (
            O => \N__62298\,
            I => \N__62197\
        );

    \I__15407\ : InMux
    port map (
            O => \N__62297\,
            I => \N__62192\
        );

    \I__15406\ : InMux
    port map (
            O => \N__62296\,
            I => \N__62192\
        );

    \I__15405\ : InMux
    port map (
            O => \N__62295\,
            I => \N__62187\
        );

    \I__15404\ : InMux
    port map (
            O => \N__62294\,
            I => \N__62187\
        );

    \I__15403\ : InMux
    port map (
            O => \N__62293\,
            I => \N__62184\
        );

    \I__15402\ : InMux
    port map (
            O => \N__62292\,
            I => \N__62179\
        );

    \I__15401\ : InMux
    port map (
            O => \N__62291\,
            I => \N__62179\
        );

    \I__15400\ : InMux
    port map (
            O => \N__62290\,
            I => \N__62176\
        );

    \I__15399\ : LocalMux
    port map (
            O => \N__62285\,
            I => \N__62171\
        );

    \I__15398\ : Span12Mux_v
    port map (
            O => \N__62276\,
            I => \N__62171\
        );

    \I__15397\ : Span4Mux_v
    port map (
            O => \N__62273\,
            I => \N__62164\
        );

    \I__15396\ : LocalMux
    port map (
            O => \N__62260\,
            I => \N__62164\
        );

    \I__15395\ : Span4Mux_v
    port map (
            O => \N__62243\,
            I => \N__62164\
        );

    \I__15394\ : InMux
    port map (
            O => \N__62242\,
            I => \N__62157\
        );

    \I__15393\ : InMux
    port map (
            O => \N__62241\,
            I => \N__62157\
        );

    \I__15392\ : InMux
    port map (
            O => \N__62240\,
            I => \N__62157\
        );

    \I__15391\ : Span4Mux_v
    port map (
            O => \N__62237\,
            I => \N__62154\
        );

    \I__15390\ : LocalMux
    port map (
            O => \N__62232\,
            I => \N__62145\
        );

    \I__15389\ : Span4Mux_h
    port map (
            O => \N__62227\,
            I => \N__62145\
        );

    \I__15388\ : Span4Mux_v
    port map (
            O => \N__62218\,
            I => \N__62145\
        );

    \I__15387\ : Span4Mux_h
    port map (
            O => \N__62215\,
            I => \N__62145\
        );

    \I__15386\ : Span4Mux_h
    port map (
            O => \N__62212\,
            I => \N__62138\
        );

    \I__15385\ : Span4Mux_h
    port map (
            O => \N__62205\,
            I => \N__62138\
        );

    \I__15384\ : Span4Mux_h
    port map (
            O => \N__62200\,
            I => \N__62138\
        );

    \I__15383\ : Odrv4
    port map (
            O => \N__62197\,
            I => comm_state_1
        );

    \I__15382\ : LocalMux
    port map (
            O => \N__62192\,
            I => comm_state_1
        );

    \I__15381\ : LocalMux
    port map (
            O => \N__62187\,
            I => comm_state_1
        );

    \I__15380\ : LocalMux
    port map (
            O => \N__62184\,
            I => comm_state_1
        );

    \I__15379\ : LocalMux
    port map (
            O => \N__62179\,
            I => comm_state_1
        );

    \I__15378\ : LocalMux
    port map (
            O => \N__62176\,
            I => comm_state_1
        );

    \I__15377\ : Odrv12
    port map (
            O => \N__62171\,
            I => comm_state_1
        );

    \I__15376\ : Odrv4
    port map (
            O => \N__62164\,
            I => comm_state_1
        );

    \I__15375\ : LocalMux
    port map (
            O => \N__62157\,
            I => comm_state_1
        );

    \I__15374\ : Odrv4
    port map (
            O => \N__62154\,
            I => comm_state_1
        );

    \I__15373\ : Odrv4
    port map (
            O => \N__62145\,
            I => comm_state_1
        );

    \I__15372\ : Odrv4
    port map (
            O => \N__62138\,
            I => comm_state_1
        );

    \I__15371\ : InMux
    port map (
            O => \N__62113\,
            I => \N__62110\
        );

    \I__15370\ : LocalMux
    port map (
            O => \N__62110\,
            I => \N__62107\
        );

    \I__15369\ : Span4Mux_h
    port map (
            O => \N__62107\,
            I => \N__62104\
        );

    \I__15368\ : Odrv4
    port map (
            O => \N__62104\,
            I => \comm_buf_0_7_N_543_3\
        );

    \I__15367\ : CascadeMux
    port map (
            O => \N__62101\,
            I => \N__62097\
        );

    \I__15366\ : CascadeMux
    port map (
            O => \N__62100\,
            I => \N__62094\
        );

    \I__15365\ : InMux
    port map (
            O => \N__62097\,
            I => \N__62087\
        );

    \I__15364\ : InMux
    port map (
            O => \N__62094\,
            I => \N__62087\
        );

    \I__15363\ : InMux
    port map (
            O => \N__62093\,
            I => \N__62083\
        );

    \I__15362\ : CascadeMux
    port map (
            O => \N__62092\,
            I => \N__62080\
        );

    \I__15361\ : LocalMux
    port map (
            O => \N__62087\,
            I => \N__62076\
        );

    \I__15360\ : InMux
    port map (
            O => \N__62086\,
            I => \N__62073\
        );

    \I__15359\ : LocalMux
    port map (
            O => \N__62083\,
            I => \N__62070\
        );

    \I__15358\ : InMux
    port map (
            O => \N__62080\,
            I => \N__62065\
        );

    \I__15357\ : InMux
    port map (
            O => \N__62079\,
            I => \N__62065\
        );

    \I__15356\ : Span4Mux_h
    port map (
            O => \N__62076\,
            I => \N__62060\
        );

    \I__15355\ : LocalMux
    port map (
            O => \N__62073\,
            I => \N__62060\
        );

    \I__15354\ : Span4Mux_v
    port map (
            O => \N__62070\,
            I => \N__62057\
        );

    \I__15353\ : LocalMux
    port map (
            O => \N__62065\,
            I => \N__62053\
        );

    \I__15352\ : Span4Mux_h
    port map (
            O => \N__62060\,
            I => \N__62050\
        );

    \I__15351\ : Span4Mux_h
    port map (
            O => \N__62057\,
            I => \N__62047\
        );

    \I__15350\ : InMux
    port map (
            O => \N__62056\,
            I => \N__62044\
        );

    \I__15349\ : Span4Mux_v
    port map (
            O => \N__62053\,
            I => \N__62041\
        );

    \I__15348\ : Span4Mux_h
    port map (
            O => \N__62050\,
            I => \N__62038\
        );

    \I__15347\ : Span4Mux_h
    port map (
            O => \N__62047\,
            I => \N__62033\
        );

    \I__15346\ : LocalMux
    port map (
            O => \N__62044\,
            I => \N__62033\
        );

    \I__15345\ : Span4Mux_h
    port map (
            O => \N__62041\,
            I => \N__62030\
        );

    \I__15344\ : Span4Mux_h
    port map (
            O => \N__62038\,
            I => \N__62025\
        );

    \I__15343\ : Span4Mux_h
    port map (
            O => \N__62033\,
            I => \N__62025\
        );

    \I__15342\ : Sp12to4
    port map (
            O => \N__62030\,
            I => \N__62022\
        );

    \I__15341\ : Span4Mux_v
    port map (
            O => \N__62025\,
            I => \N__62019\
        );

    \I__15340\ : Odrv12
    port map (
            O => \N__62022\,
            I => comm_buf_0_3
        );

    \I__15339\ : Odrv4
    port map (
            O => \N__62019\,
            I => comm_buf_0_3
        );

    \I__15338\ : ClkMux
    port map (
            O => \N__62014\,
            I => \N__61441\
        );

    \I__15337\ : ClkMux
    port map (
            O => \N__62013\,
            I => \N__61441\
        );

    \I__15336\ : ClkMux
    port map (
            O => \N__62012\,
            I => \N__61441\
        );

    \I__15335\ : ClkMux
    port map (
            O => \N__62011\,
            I => \N__61441\
        );

    \I__15334\ : ClkMux
    port map (
            O => \N__62010\,
            I => \N__61441\
        );

    \I__15333\ : ClkMux
    port map (
            O => \N__62009\,
            I => \N__61441\
        );

    \I__15332\ : ClkMux
    port map (
            O => \N__62008\,
            I => \N__61441\
        );

    \I__15331\ : ClkMux
    port map (
            O => \N__62007\,
            I => \N__61441\
        );

    \I__15330\ : ClkMux
    port map (
            O => \N__62006\,
            I => \N__61441\
        );

    \I__15329\ : ClkMux
    port map (
            O => \N__62005\,
            I => \N__61441\
        );

    \I__15328\ : ClkMux
    port map (
            O => \N__62004\,
            I => \N__61441\
        );

    \I__15327\ : ClkMux
    port map (
            O => \N__62003\,
            I => \N__61441\
        );

    \I__15326\ : ClkMux
    port map (
            O => \N__62002\,
            I => \N__61441\
        );

    \I__15325\ : ClkMux
    port map (
            O => \N__62001\,
            I => \N__61441\
        );

    \I__15324\ : ClkMux
    port map (
            O => \N__62000\,
            I => \N__61441\
        );

    \I__15323\ : ClkMux
    port map (
            O => \N__61999\,
            I => \N__61441\
        );

    \I__15322\ : ClkMux
    port map (
            O => \N__61998\,
            I => \N__61441\
        );

    \I__15321\ : ClkMux
    port map (
            O => \N__61997\,
            I => \N__61441\
        );

    \I__15320\ : ClkMux
    port map (
            O => \N__61996\,
            I => \N__61441\
        );

    \I__15319\ : ClkMux
    port map (
            O => \N__61995\,
            I => \N__61441\
        );

    \I__15318\ : ClkMux
    port map (
            O => \N__61994\,
            I => \N__61441\
        );

    \I__15317\ : ClkMux
    port map (
            O => \N__61993\,
            I => \N__61441\
        );

    \I__15316\ : ClkMux
    port map (
            O => \N__61992\,
            I => \N__61441\
        );

    \I__15315\ : ClkMux
    port map (
            O => \N__61991\,
            I => \N__61441\
        );

    \I__15314\ : ClkMux
    port map (
            O => \N__61990\,
            I => \N__61441\
        );

    \I__15313\ : ClkMux
    port map (
            O => \N__61989\,
            I => \N__61441\
        );

    \I__15312\ : ClkMux
    port map (
            O => \N__61988\,
            I => \N__61441\
        );

    \I__15311\ : ClkMux
    port map (
            O => \N__61987\,
            I => \N__61441\
        );

    \I__15310\ : ClkMux
    port map (
            O => \N__61986\,
            I => \N__61441\
        );

    \I__15309\ : ClkMux
    port map (
            O => \N__61985\,
            I => \N__61441\
        );

    \I__15308\ : ClkMux
    port map (
            O => \N__61984\,
            I => \N__61441\
        );

    \I__15307\ : ClkMux
    port map (
            O => \N__61983\,
            I => \N__61441\
        );

    \I__15306\ : ClkMux
    port map (
            O => \N__61982\,
            I => \N__61441\
        );

    \I__15305\ : ClkMux
    port map (
            O => \N__61981\,
            I => \N__61441\
        );

    \I__15304\ : ClkMux
    port map (
            O => \N__61980\,
            I => \N__61441\
        );

    \I__15303\ : ClkMux
    port map (
            O => \N__61979\,
            I => \N__61441\
        );

    \I__15302\ : ClkMux
    port map (
            O => \N__61978\,
            I => \N__61441\
        );

    \I__15301\ : ClkMux
    port map (
            O => \N__61977\,
            I => \N__61441\
        );

    \I__15300\ : ClkMux
    port map (
            O => \N__61976\,
            I => \N__61441\
        );

    \I__15299\ : ClkMux
    port map (
            O => \N__61975\,
            I => \N__61441\
        );

    \I__15298\ : ClkMux
    port map (
            O => \N__61974\,
            I => \N__61441\
        );

    \I__15297\ : ClkMux
    port map (
            O => \N__61973\,
            I => \N__61441\
        );

    \I__15296\ : ClkMux
    port map (
            O => \N__61972\,
            I => \N__61441\
        );

    \I__15295\ : ClkMux
    port map (
            O => \N__61971\,
            I => \N__61441\
        );

    \I__15294\ : ClkMux
    port map (
            O => \N__61970\,
            I => \N__61441\
        );

    \I__15293\ : ClkMux
    port map (
            O => \N__61969\,
            I => \N__61441\
        );

    \I__15292\ : ClkMux
    port map (
            O => \N__61968\,
            I => \N__61441\
        );

    \I__15291\ : ClkMux
    port map (
            O => \N__61967\,
            I => \N__61441\
        );

    \I__15290\ : ClkMux
    port map (
            O => \N__61966\,
            I => \N__61441\
        );

    \I__15289\ : ClkMux
    port map (
            O => \N__61965\,
            I => \N__61441\
        );

    \I__15288\ : ClkMux
    port map (
            O => \N__61964\,
            I => \N__61441\
        );

    \I__15287\ : ClkMux
    port map (
            O => \N__61963\,
            I => \N__61441\
        );

    \I__15286\ : ClkMux
    port map (
            O => \N__61962\,
            I => \N__61441\
        );

    \I__15285\ : ClkMux
    port map (
            O => \N__61961\,
            I => \N__61441\
        );

    \I__15284\ : ClkMux
    port map (
            O => \N__61960\,
            I => \N__61441\
        );

    \I__15283\ : ClkMux
    port map (
            O => \N__61959\,
            I => \N__61441\
        );

    \I__15282\ : ClkMux
    port map (
            O => \N__61958\,
            I => \N__61441\
        );

    \I__15281\ : ClkMux
    port map (
            O => \N__61957\,
            I => \N__61441\
        );

    \I__15280\ : ClkMux
    port map (
            O => \N__61956\,
            I => \N__61441\
        );

    \I__15279\ : ClkMux
    port map (
            O => \N__61955\,
            I => \N__61441\
        );

    \I__15278\ : ClkMux
    port map (
            O => \N__61954\,
            I => \N__61441\
        );

    \I__15277\ : ClkMux
    port map (
            O => \N__61953\,
            I => \N__61441\
        );

    \I__15276\ : ClkMux
    port map (
            O => \N__61952\,
            I => \N__61441\
        );

    \I__15275\ : ClkMux
    port map (
            O => \N__61951\,
            I => \N__61441\
        );

    \I__15274\ : ClkMux
    port map (
            O => \N__61950\,
            I => \N__61441\
        );

    \I__15273\ : ClkMux
    port map (
            O => \N__61949\,
            I => \N__61441\
        );

    \I__15272\ : ClkMux
    port map (
            O => \N__61948\,
            I => \N__61441\
        );

    \I__15271\ : ClkMux
    port map (
            O => \N__61947\,
            I => \N__61441\
        );

    \I__15270\ : ClkMux
    port map (
            O => \N__61946\,
            I => \N__61441\
        );

    \I__15269\ : ClkMux
    port map (
            O => \N__61945\,
            I => \N__61441\
        );

    \I__15268\ : ClkMux
    port map (
            O => \N__61944\,
            I => \N__61441\
        );

    \I__15267\ : ClkMux
    port map (
            O => \N__61943\,
            I => \N__61441\
        );

    \I__15266\ : ClkMux
    port map (
            O => \N__61942\,
            I => \N__61441\
        );

    \I__15265\ : ClkMux
    port map (
            O => \N__61941\,
            I => \N__61441\
        );

    \I__15264\ : ClkMux
    port map (
            O => \N__61940\,
            I => \N__61441\
        );

    \I__15263\ : ClkMux
    port map (
            O => \N__61939\,
            I => \N__61441\
        );

    \I__15262\ : ClkMux
    port map (
            O => \N__61938\,
            I => \N__61441\
        );

    \I__15261\ : ClkMux
    port map (
            O => \N__61937\,
            I => \N__61441\
        );

    \I__15260\ : ClkMux
    port map (
            O => \N__61936\,
            I => \N__61441\
        );

    \I__15259\ : ClkMux
    port map (
            O => \N__61935\,
            I => \N__61441\
        );

    \I__15258\ : ClkMux
    port map (
            O => \N__61934\,
            I => \N__61441\
        );

    \I__15257\ : ClkMux
    port map (
            O => \N__61933\,
            I => \N__61441\
        );

    \I__15256\ : ClkMux
    port map (
            O => \N__61932\,
            I => \N__61441\
        );

    \I__15255\ : ClkMux
    port map (
            O => \N__61931\,
            I => \N__61441\
        );

    \I__15254\ : ClkMux
    port map (
            O => \N__61930\,
            I => \N__61441\
        );

    \I__15253\ : ClkMux
    port map (
            O => \N__61929\,
            I => \N__61441\
        );

    \I__15252\ : ClkMux
    port map (
            O => \N__61928\,
            I => \N__61441\
        );

    \I__15251\ : ClkMux
    port map (
            O => \N__61927\,
            I => \N__61441\
        );

    \I__15250\ : ClkMux
    port map (
            O => \N__61926\,
            I => \N__61441\
        );

    \I__15249\ : ClkMux
    port map (
            O => \N__61925\,
            I => \N__61441\
        );

    \I__15248\ : ClkMux
    port map (
            O => \N__61924\,
            I => \N__61441\
        );

    \I__15247\ : ClkMux
    port map (
            O => \N__61923\,
            I => \N__61441\
        );

    \I__15246\ : ClkMux
    port map (
            O => \N__61922\,
            I => \N__61441\
        );

    \I__15245\ : ClkMux
    port map (
            O => \N__61921\,
            I => \N__61441\
        );

    \I__15244\ : ClkMux
    port map (
            O => \N__61920\,
            I => \N__61441\
        );

    \I__15243\ : ClkMux
    port map (
            O => \N__61919\,
            I => \N__61441\
        );

    \I__15242\ : ClkMux
    port map (
            O => \N__61918\,
            I => \N__61441\
        );

    \I__15241\ : ClkMux
    port map (
            O => \N__61917\,
            I => \N__61441\
        );

    \I__15240\ : ClkMux
    port map (
            O => \N__61916\,
            I => \N__61441\
        );

    \I__15239\ : ClkMux
    port map (
            O => \N__61915\,
            I => \N__61441\
        );

    \I__15238\ : ClkMux
    port map (
            O => \N__61914\,
            I => \N__61441\
        );

    \I__15237\ : ClkMux
    port map (
            O => \N__61913\,
            I => \N__61441\
        );

    \I__15236\ : ClkMux
    port map (
            O => \N__61912\,
            I => \N__61441\
        );

    \I__15235\ : ClkMux
    port map (
            O => \N__61911\,
            I => \N__61441\
        );

    \I__15234\ : ClkMux
    port map (
            O => \N__61910\,
            I => \N__61441\
        );

    \I__15233\ : ClkMux
    port map (
            O => \N__61909\,
            I => \N__61441\
        );

    \I__15232\ : ClkMux
    port map (
            O => \N__61908\,
            I => \N__61441\
        );

    \I__15231\ : ClkMux
    port map (
            O => \N__61907\,
            I => \N__61441\
        );

    \I__15230\ : ClkMux
    port map (
            O => \N__61906\,
            I => \N__61441\
        );

    \I__15229\ : ClkMux
    port map (
            O => \N__61905\,
            I => \N__61441\
        );

    \I__15228\ : ClkMux
    port map (
            O => \N__61904\,
            I => \N__61441\
        );

    \I__15227\ : ClkMux
    port map (
            O => \N__61903\,
            I => \N__61441\
        );

    \I__15226\ : ClkMux
    port map (
            O => \N__61902\,
            I => \N__61441\
        );

    \I__15225\ : ClkMux
    port map (
            O => \N__61901\,
            I => \N__61441\
        );

    \I__15224\ : ClkMux
    port map (
            O => \N__61900\,
            I => \N__61441\
        );

    \I__15223\ : ClkMux
    port map (
            O => \N__61899\,
            I => \N__61441\
        );

    \I__15222\ : ClkMux
    port map (
            O => \N__61898\,
            I => \N__61441\
        );

    \I__15221\ : ClkMux
    port map (
            O => \N__61897\,
            I => \N__61441\
        );

    \I__15220\ : ClkMux
    port map (
            O => \N__61896\,
            I => \N__61441\
        );

    \I__15219\ : ClkMux
    port map (
            O => \N__61895\,
            I => \N__61441\
        );

    \I__15218\ : ClkMux
    port map (
            O => \N__61894\,
            I => \N__61441\
        );

    \I__15217\ : ClkMux
    port map (
            O => \N__61893\,
            I => \N__61441\
        );

    \I__15216\ : ClkMux
    port map (
            O => \N__61892\,
            I => \N__61441\
        );

    \I__15215\ : ClkMux
    port map (
            O => \N__61891\,
            I => \N__61441\
        );

    \I__15214\ : ClkMux
    port map (
            O => \N__61890\,
            I => \N__61441\
        );

    \I__15213\ : ClkMux
    port map (
            O => \N__61889\,
            I => \N__61441\
        );

    \I__15212\ : ClkMux
    port map (
            O => \N__61888\,
            I => \N__61441\
        );

    \I__15211\ : ClkMux
    port map (
            O => \N__61887\,
            I => \N__61441\
        );

    \I__15210\ : ClkMux
    port map (
            O => \N__61886\,
            I => \N__61441\
        );

    \I__15209\ : ClkMux
    port map (
            O => \N__61885\,
            I => \N__61441\
        );

    \I__15208\ : ClkMux
    port map (
            O => \N__61884\,
            I => \N__61441\
        );

    \I__15207\ : ClkMux
    port map (
            O => \N__61883\,
            I => \N__61441\
        );

    \I__15206\ : ClkMux
    port map (
            O => \N__61882\,
            I => \N__61441\
        );

    \I__15205\ : ClkMux
    port map (
            O => \N__61881\,
            I => \N__61441\
        );

    \I__15204\ : ClkMux
    port map (
            O => \N__61880\,
            I => \N__61441\
        );

    \I__15203\ : ClkMux
    port map (
            O => \N__61879\,
            I => \N__61441\
        );

    \I__15202\ : ClkMux
    port map (
            O => \N__61878\,
            I => \N__61441\
        );

    \I__15201\ : ClkMux
    port map (
            O => \N__61877\,
            I => \N__61441\
        );

    \I__15200\ : ClkMux
    port map (
            O => \N__61876\,
            I => \N__61441\
        );

    \I__15199\ : ClkMux
    port map (
            O => \N__61875\,
            I => \N__61441\
        );

    \I__15198\ : ClkMux
    port map (
            O => \N__61874\,
            I => \N__61441\
        );

    \I__15197\ : ClkMux
    port map (
            O => \N__61873\,
            I => \N__61441\
        );

    \I__15196\ : ClkMux
    port map (
            O => \N__61872\,
            I => \N__61441\
        );

    \I__15195\ : ClkMux
    port map (
            O => \N__61871\,
            I => \N__61441\
        );

    \I__15194\ : ClkMux
    port map (
            O => \N__61870\,
            I => \N__61441\
        );

    \I__15193\ : ClkMux
    port map (
            O => \N__61869\,
            I => \N__61441\
        );

    \I__15192\ : ClkMux
    port map (
            O => \N__61868\,
            I => \N__61441\
        );

    \I__15191\ : ClkMux
    port map (
            O => \N__61867\,
            I => \N__61441\
        );

    \I__15190\ : ClkMux
    port map (
            O => \N__61866\,
            I => \N__61441\
        );

    \I__15189\ : ClkMux
    port map (
            O => \N__61865\,
            I => \N__61441\
        );

    \I__15188\ : ClkMux
    port map (
            O => \N__61864\,
            I => \N__61441\
        );

    \I__15187\ : ClkMux
    port map (
            O => \N__61863\,
            I => \N__61441\
        );

    \I__15186\ : ClkMux
    port map (
            O => \N__61862\,
            I => \N__61441\
        );

    \I__15185\ : ClkMux
    port map (
            O => \N__61861\,
            I => \N__61441\
        );

    \I__15184\ : ClkMux
    port map (
            O => \N__61860\,
            I => \N__61441\
        );

    \I__15183\ : ClkMux
    port map (
            O => \N__61859\,
            I => \N__61441\
        );

    \I__15182\ : ClkMux
    port map (
            O => \N__61858\,
            I => \N__61441\
        );

    \I__15181\ : ClkMux
    port map (
            O => \N__61857\,
            I => \N__61441\
        );

    \I__15180\ : ClkMux
    port map (
            O => \N__61856\,
            I => \N__61441\
        );

    \I__15179\ : ClkMux
    port map (
            O => \N__61855\,
            I => \N__61441\
        );

    \I__15178\ : ClkMux
    port map (
            O => \N__61854\,
            I => \N__61441\
        );

    \I__15177\ : ClkMux
    port map (
            O => \N__61853\,
            I => \N__61441\
        );

    \I__15176\ : ClkMux
    port map (
            O => \N__61852\,
            I => \N__61441\
        );

    \I__15175\ : ClkMux
    port map (
            O => \N__61851\,
            I => \N__61441\
        );

    \I__15174\ : ClkMux
    port map (
            O => \N__61850\,
            I => \N__61441\
        );

    \I__15173\ : ClkMux
    port map (
            O => \N__61849\,
            I => \N__61441\
        );

    \I__15172\ : ClkMux
    port map (
            O => \N__61848\,
            I => \N__61441\
        );

    \I__15171\ : ClkMux
    port map (
            O => \N__61847\,
            I => \N__61441\
        );

    \I__15170\ : ClkMux
    port map (
            O => \N__61846\,
            I => \N__61441\
        );

    \I__15169\ : ClkMux
    port map (
            O => \N__61845\,
            I => \N__61441\
        );

    \I__15168\ : ClkMux
    port map (
            O => \N__61844\,
            I => \N__61441\
        );

    \I__15167\ : ClkMux
    port map (
            O => \N__61843\,
            I => \N__61441\
        );

    \I__15166\ : ClkMux
    port map (
            O => \N__61842\,
            I => \N__61441\
        );

    \I__15165\ : ClkMux
    port map (
            O => \N__61841\,
            I => \N__61441\
        );

    \I__15164\ : ClkMux
    port map (
            O => \N__61840\,
            I => \N__61441\
        );

    \I__15163\ : ClkMux
    port map (
            O => \N__61839\,
            I => \N__61441\
        );

    \I__15162\ : ClkMux
    port map (
            O => \N__61838\,
            I => \N__61441\
        );

    \I__15161\ : ClkMux
    port map (
            O => \N__61837\,
            I => \N__61441\
        );

    \I__15160\ : ClkMux
    port map (
            O => \N__61836\,
            I => \N__61441\
        );

    \I__15159\ : ClkMux
    port map (
            O => \N__61835\,
            I => \N__61441\
        );

    \I__15158\ : ClkMux
    port map (
            O => \N__61834\,
            I => \N__61441\
        );

    \I__15157\ : ClkMux
    port map (
            O => \N__61833\,
            I => \N__61441\
        );

    \I__15156\ : ClkMux
    port map (
            O => \N__61832\,
            I => \N__61441\
        );

    \I__15155\ : ClkMux
    port map (
            O => \N__61831\,
            I => \N__61441\
        );

    \I__15154\ : ClkMux
    port map (
            O => \N__61830\,
            I => \N__61441\
        );

    \I__15153\ : ClkMux
    port map (
            O => \N__61829\,
            I => \N__61441\
        );

    \I__15152\ : ClkMux
    port map (
            O => \N__61828\,
            I => \N__61441\
        );

    \I__15151\ : ClkMux
    port map (
            O => \N__61827\,
            I => \N__61441\
        );

    \I__15150\ : ClkMux
    port map (
            O => \N__61826\,
            I => \N__61441\
        );

    \I__15149\ : ClkMux
    port map (
            O => \N__61825\,
            I => \N__61441\
        );

    \I__15148\ : ClkMux
    port map (
            O => \N__61824\,
            I => \N__61441\
        );

    \I__15147\ : GlobalMux
    port map (
            O => \N__61441\,
            I => \clk_32MHz\
        );

    \I__15146\ : CEMux
    port map (
            O => \N__61438\,
            I => \N__61434\
        );

    \I__15145\ : CEMux
    port map (
            O => \N__61437\,
            I => \N__61431\
        );

    \I__15144\ : LocalMux
    port map (
            O => \N__61434\,
            I => \N__61428\
        );

    \I__15143\ : LocalMux
    port map (
            O => \N__61431\,
            I => \N__61425\
        );

    \I__15142\ : Span4Mux_h
    port map (
            O => \N__61428\,
            I => \N__61420\
        );

    \I__15141\ : Span4Mux_h
    port map (
            O => \N__61425\,
            I => \N__61420\
        );

    \I__15140\ : Odrv4
    port map (
            O => \N__61420\,
            I => n12677
        );

    \I__15139\ : CascadeMux
    port map (
            O => \N__61417\,
            I => \n30_adj_1793_cascade_\
        );

    \I__15138\ : CascadeMux
    port map (
            O => \N__61414\,
            I => \N__61402\
        );

    \I__15137\ : CascadeMux
    port map (
            O => \N__61413\,
            I => \N__61391\
        );

    \I__15136\ : InMux
    port map (
            O => \N__61412\,
            I => \N__61387\
        );

    \I__15135\ : InMux
    port map (
            O => \N__61411\,
            I => \N__61384\
        );

    \I__15134\ : InMux
    port map (
            O => \N__61410\,
            I => \N__61376\
        );

    \I__15133\ : InMux
    port map (
            O => \N__61409\,
            I => \N__61370\
        );

    \I__15132\ : InMux
    port map (
            O => \N__61408\,
            I => \N__61367\
        );

    \I__15131\ : InMux
    port map (
            O => \N__61407\,
            I => \N__61364\
        );

    \I__15130\ : InMux
    port map (
            O => \N__61406\,
            I => \N__61359\
        );

    \I__15129\ : InMux
    port map (
            O => \N__61405\,
            I => \N__61356\
        );

    \I__15128\ : InMux
    port map (
            O => \N__61402\,
            I => \N__61353\
        );

    \I__15127\ : InMux
    port map (
            O => \N__61401\,
            I => \N__61349\
        );

    \I__15126\ : InMux
    port map (
            O => \N__61400\,
            I => \N__61344\
        );

    \I__15125\ : InMux
    port map (
            O => \N__61399\,
            I => \N__61339\
        );

    \I__15124\ : InMux
    port map (
            O => \N__61398\,
            I => \N__61339\
        );

    \I__15123\ : InMux
    port map (
            O => \N__61397\,
            I => \N__61336\
        );

    \I__15122\ : InMux
    port map (
            O => \N__61396\,
            I => \N__61333\
        );

    \I__15121\ : InMux
    port map (
            O => \N__61395\,
            I => \N__61330\
        );

    \I__15120\ : InMux
    port map (
            O => \N__61394\,
            I => \N__61327\
        );

    \I__15119\ : InMux
    port map (
            O => \N__61391\,
            I => \N__61322\
        );

    \I__15118\ : InMux
    port map (
            O => \N__61390\,
            I => \N__61322\
        );

    \I__15117\ : LocalMux
    port map (
            O => \N__61387\,
            I => \N__61319\
        );

    \I__15116\ : LocalMux
    port map (
            O => \N__61384\,
            I => \N__61316\
        );

    \I__15115\ : InMux
    port map (
            O => \N__61383\,
            I => \N__61313\
        );

    \I__15114\ : InMux
    port map (
            O => \N__61382\,
            I => \N__61310\
        );

    \I__15113\ : InMux
    port map (
            O => \N__61381\,
            I => \N__61307\
        );

    \I__15112\ : InMux
    port map (
            O => \N__61380\,
            I => \N__61304\
        );

    \I__15111\ : InMux
    port map (
            O => \N__61379\,
            I => \N__61301\
        );

    \I__15110\ : LocalMux
    port map (
            O => \N__61376\,
            I => \N__61297\
        );

    \I__15109\ : InMux
    port map (
            O => \N__61375\,
            I => \N__61292\
        );

    \I__15108\ : InMux
    port map (
            O => \N__61374\,
            I => \N__61292\
        );

    \I__15107\ : InMux
    port map (
            O => \N__61373\,
            I => \N__61288\
        );

    \I__15106\ : LocalMux
    port map (
            O => \N__61370\,
            I => \N__61281\
        );

    \I__15105\ : LocalMux
    port map (
            O => \N__61367\,
            I => \N__61281\
        );

    \I__15104\ : LocalMux
    port map (
            O => \N__61364\,
            I => \N__61281\
        );

    \I__15103\ : InMux
    port map (
            O => \N__61363\,
            I => \N__61276\
        );

    \I__15102\ : InMux
    port map (
            O => \N__61362\,
            I => \N__61276\
        );

    \I__15101\ : LocalMux
    port map (
            O => \N__61359\,
            I => \N__61269\
        );

    \I__15100\ : LocalMux
    port map (
            O => \N__61356\,
            I => \N__61269\
        );

    \I__15099\ : LocalMux
    port map (
            O => \N__61353\,
            I => \N__61269\
        );

    \I__15098\ : InMux
    port map (
            O => \N__61352\,
            I => \N__61264\
        );

    \I__15097\ : LocalMux
    port map (
            O => \N__61349\,
            I => \N__61261\
        );

    \I__15096\ : InMux
    port map (
            O => \N__61348\,
            I => \N__61255\
        );

    \I__15095\ : InMux
    port map (
            O => \N__61347\,
            I => \N__61255\
        );

    \I__15094\ : LocalMux
    port map (
            O => \N__61344\,
            I => \N__61248\
        );

    \I__15093\ : LocalMux
    port map (
            O => \N__61339\,
            I => \N__61248\
        );

    \I__15092\ : LocalMux
    port map (
            O => \N__61336\,
            I => \N__61245\
        );

    \I__15091\ : LocalMux
    port map (
            O => \N__61333\,
            I => \N__61242\
        );

    \I__15090\ : LocalMux
    port map (
            O => \N__61330\,
            I => \N__61233\
        );

    \I__15089\ : LocalMux
    port map (
            O => \N__61327\,
            I => \N__61233\
        );

    \I__15088\ : LocalMux
    port map (
            O => \N__61322\,
            I => \N__61233\
        );

    \I__15087\ : Span4Mux_v
    port map (
            O => \N__61319\,
            I => \N__61233\
        );

    \I__15086\ : Span4Mux_h
    port map (
            O => \N__61316\,
            I => \N__61226\
        );

    \I__15085\ : LocalMux
    port map (
            O => \N__61313\,
            I => \N__61226\
        );

    \I__15084\ : LocalMux
    port map (
            O => \N__61310\,
            I => \N__61223\
        );

    \I__15083\ : LocalMux
    port map (
            O => \N__61307\,
            I => \N__61218\
        );

    \I__15082\ : LocalMux
    port map (
            O => \N__61304\,
            I => \N__61218\
        );

    \I__15081\ : LocalMux
    port map (
            O => \N__61301\,
            I => \N__61215\
        );

    \I__15080\ : InMux
    port map (
            O => \N__61300\,
            I => \N__61212\
        );

    \I__15079\ : Span4Mux_v
    port map (
            O => \N__61297\,
            I => \N__61207\
        );

    \I__15078\ : LocalMux
    port map (
            O => \N__61292\,
            I => \N__61207\
        );

    \I__15077\ : InMux
    port map (
            O => \N__61291\,
            I => \N__61204\
        );

    \I__15076\ : LocalMux
    port map (
            O => \N__61288\,
            I => \N__61201\
        );

    \I__15075\ : Span4Mux_v
    port map (
            O => \N__61281\,
            I => \N__61194\
        );

    \I__15074\ : LocalMux
    port map (
            O => \N__61276\,
            I => \N__61194\
        );

    \I__15073\ : Span4Mux_h
    port map (
            O => \N__61269\,
            I => \N__61194\
        );

    \I__15072\ : InMux
    port map (
            O => \N__61268\,
            I => \N__61189\
        );

    \I__15071\ : InMux
    port map (
            O => \N__61267\,
            I => \N__61189\
        );

    \I__15070\ : LocalMux
    port map (
            O => \N__61264\,
            I => \N__61184\
        );

    \I__15069\ : Span4Mux_h
    port map (
            O => \N__61261\,
            I => \N__61184\
        );

    \I__15068\ : CascadeMux
    port map (
            O => \N__61260\,
            I => \N__61179\
        );

    \I__15067\ : LocalMux
    port map (
            O => \N__61255\,
            I => \N__61175\
        );

    \I__15066\ : InMux
    port map (
            O => \N__61254\,
            I => \N__61172\
        );

    \I__15065\ : InMux
    port map (
            O => \N__61253\,
            I => \N__61169\
        );

    \I__15064\ : Span4Mux_v
    port map (
            O => \N__61248\,
            I => \N__61160\
        );

    \I__15063\ : Span4Mux_v
    port map (
            O => \N__61245\,
            I => \N__61160\
        );

    \I__15062\ : Span4Mux_v
    port map (
            O => \N__61242\,
            I => \N__61160\
        );

    \I__15061\ : Span4Mux_h
    port map (
            O => \N__61233\,
            I => \N__61160\
        );

    \I__15060\ : InMux
    port map (
            O => \N__61232\,
            I => \N__61157\
        );

    \I__15059\ : InMux
    port map (
            O => \N__61231\,
            I => \N__61154\
        );

    \I__15058\ : Span4Mux_v
    port map (
            O => \N__61226\,
            I => \N__61141\
        );

    \I__15057\ : Span4Mux_v
    port map (
            O => \N__61223\,
            I => \N__61141\
        );

    \I__15056\ : Span4Mux_v
    port map (
            O => \N__61218\,
            I => \N__61141\
        );

    \I__15055\ : Span4Mux_h
    port map (
            O => \N__61215\,
            I => \N__61141\
        );

    \I__15054\ : LocalMux
    port map (
            O => \N__61212\,
            I => \N__61141\
        );

    \I__15053\ : Span4Mux_h
    port map (
            O => \N__61207\,
            I => \N__61141\
        );

    \I__15052\ : LocalMux
    port map (
            O => \N__61204\,
            I => \N__61130\
        );

    \I__15051\ : Span4Mux_v
    port map (
            O => \N__61201\,
            I => \N__61130\
        );

    \I__15050\ : Span4Mux_h
    port map (
            O => \N__61194\,
            I => \N__61130\
        );

    \I__15049\ : LocalMux
    port map (
            O => \N__61189\,
            I => \N__61130\
        );

    \I__15048\ : Span4Mux_h
    port map (
            O => \N__61184\,
            I => \N__61130\
        );

    \I__15047\ : InMux
    port map (
            O => \N__61183\,
            I => \N__61121\
        );

    \I__15046\ : InMux
    port map (
            O => \N__61182\,
            I => \N__61121\
        );

    \I__15045\ : InMux
    port map (
            O => \N__61179\,
            I => \N__61121\
        );

    \I__15044\ : InMux
    port map (
            O => \N__61178\,
            I => \N__61121\
        );

    \I__15043\ : Odrv12
    port map (
            O => \N__61175\,
            I => comm_cmd_6
        );

    \I__15042\ : LocalMux
    port map (
            O => \N__61172\,
            I => comm_cmd_6
        );

    \I__15041\ : LocalMux
    port map (
            O => \N__61169\,
            I => comm_cmd_6
        );

    \I__15040\ : Odrv4
    port map (
            O => \N__61160\,
            I => comm_cmd_6
        );

    \I__15039\ : LocalMux
    port map (
            O => \N__61157\,
            I => comm_cmd_6
        );

    \I__15038\ : LocalMux
    port map (
            O => \N__61154\,
            I => comm_cmd_6
        );

    \I__15037\ : Odrv4
    port map (
            O => \N__61141\,
            I => comm_cmd_6
        );

    \I__15036\ : Odrv4
    port map (
            O => \N__61130\,
            I => comm_cmd_6
        );

    \I__15035\ : LocalMux
    port map (
            O => \N__61121\,
            I => comm_cmd_6
        );

    \I__15034\ : CascadeMux
    port map (
            O => \N__61102\,
            I => \N__61099\
        );

    \I__15033\ : InMux
    port map (
            O => \N__61099\,
            I => \N__61096\
        );

    \I__15032\ : LocalMux
    port map (
            O => \N__61096\,
            I => \N__61092\
        );

    \I__15031\ : CascadeMux
    port map (
            O => \N__61095\,
            I => \N__61089\
        );

    \I__15030\ : Span4Mux_v
    port map (
            O => \N__61092\,
            I => \N__61086\
        );

    \I__15029\ : InMux
    port map (
            O => \N__61089\,
            I => \N__61083\
        );

    \I__15028\ : Span4Mux_h
    port map (
            O => \N__61086\,
            I => \N__61080\
        );

    \I__15027\ : LocalMux
    port map (
            O => \N__61083\,
            I => data_idxvec_13
        );

    \I__15026\ : Odrv4
    port map (
            O => \N__61080\,
            I => data_idxvec_13
        );

    \I__15025\ : InMux
    port map (
            O => \N__61075\,
            I => \N__61072\
        );

    \I__15024\ : LocalMux
    port map (
            O => \N__61072\,
            I => \N__61069\
        );

    \I__15023\ : Span4Mux_v
    port map (
            O => \N__61069\,
            I => \N__61066\
        );

    \I__15022\ : Span4Mux_v
    port map (
            O => \N__61066\,
            I => \N__61063\
        );

    \I__15021\ : Odrv4
    port map (
            O => \N__61063\,
            I => buf_data_iac_21
        );

    \I__15020\ : CascadeMux
    port map (
            O => \N__61060\,
            I => \n28_adj_1775_cascade_\
        );

    \I__15019\ : CascadeMux
    port map (
            O => \N__61057\,
            I => \N__61048\
        );

    \I__15018\ : InMux
    port map (
            O => \N__61056\,
            I => \N__61045\
        );

    \I__15017\ : InMux
    port map (
            O => \N__61055\,
            I => \N__61042\
        );

    \I__15016\ : InMux
    port map (
            O => \N__61054\,
            I => \N__61037\
        );

    \I__15015\ : InMux
    port map (
            O => \N__61053\,
            I => \N__61037\
        );

    \I__15014\ : InMux
    port map (
            O => \N__61052\,
            I => \N__61029\
        );

    \I__15013\ : InMux
    port map (
            O => \N__61051\,
            I => \N__61026\
        );

    \I__15012\ : InMux
    port map (
            O => \N__61048\,
            I => \N__61014\
        );

    \I__15011\ : LocalMux
    port map (
            O => \N__61045\,
            I => \N__61010\
        );

    \I__15010\ : LocalMux
    port map (
            O => \N__61042\,
            I => \N__61007\
        );

    \I__15009\ : LocalMux
    port map (
            O => \N__61037\,
            I => \N__61004\
        );

    \I__15008\ : InMux
    port map (
            O => \N__61036\,
            I => \N__60995\
        );

    \I__15007\ : InMux
    port map (
            O => \N__61035\,
            I => \N__60995\
        );

    \I__15006\ : InMux
    port map (
            O => \N__61034\,
            I => \N__60995\
        );

    \I__15005\ : InMux
    port map (
            O => \N__61033\,
            I => \N__60995\
        );

    \I__15004\ : InMux
    port map (
            O => \N__61032\,
            I => \N__60986\
        );

    \I__15003\ : LocalMux
    port map (
            O => \N__61029\,
            I => \N__60981\
        );

    \I__15002\ : LocalMux
    port map (
            O => \N__61026\,
            I => \N__60981\
        );

    \I__15001\ : InMux
    port map (
            O => \N__61025\,
            I => \N__60970\
        );

    \I__15000\ : InMux
    port map (
            O => \N__61024\,
            I => \N__60970\
        );

    \I__14999\ : InMux
    port map (
            O => \N__61023\,
            I => \N__60963\
        );

    \I__14998\ : InMux
    port map (
            O => \N__61022\,
            I => \N__60963\
        );

    \I__14997\ : InMux
    port map (
            O => \N__61021\,
            I => \N__60963\
        );

    \I__14996\ : InMux
    port map (
            O => \N__61020\,
            I => \N__60958\
        );

    \I__14995\ : InMux
    port map (
            O => \N__61019\,
            I => \N__60958\
        );

    \I__14994\ : CascadeMux
    port map (
            O => \N__61018\,
            I => \N__60949\
        );

    \I__14993\ : InMux
    port map (
            O => \N__61017\,
            I => \N__60945\
        );

    \I__14992\ : LocalMux
    port map (
            O => \N__61014\,
            I => \N__60942\
        );

    \I__14991\ : InMux
    port map (
            O => \N__61013\,
            I => \N__60939\
        );

    \I__14990\ : Span4Mux_v
    port map (
            O => \N__61010\,
            I => \N__60932\
        );

    \I__14989\ : Span4Mux_v
    port map (
            O => \N__61007\,
            I => \N__60932\
        );

    \I__14988\ : Span4Mux_h
    port map (
            O => \N__61004\,
            I => \N__60932\
        );

    \I__14987\ : LocalMux
    port map (
            O => \N__60995\,
            I => \N__60929\
        );

    \I__14986\ : InMux
    port map (
            O => \N__60994\,
            I => \N__60926\
        );

    \I__14985\ : InMux
    port map (
            O => \N__60993\,
            I => \N__60921\
        );

    \I__14984\ : InMux
    port map (
            O => \N__60992\,
            I => \N__60921\
        );

    \I__14983\ : InMux
    port map (
            O => \N__60991\,
            I => \N__60918\
        );

    \I__14982\ : InMux
    port map (
            O => \N__60990\,
            I => \N__60915\
        );

    \I__14981\ : InMux
    port map (
            O => \N__60989\,
            I => \N__60912\
        );

    \I__14980\ : LocalMux
    port map (
            O => \N__60986\,
            I => \N__60909\
        );

    \I__14979\ : Span4Mux_v
    port map (
            O => \N__60981\,
            I => \N__60906\
        );

    \I__14978\ : InMux
    port map (
            O => \N__60980\,
            I => \N__60903\
        );

    \I__14977\ : InMux
    port map (
            O => \N__60979\,
            I => \N__60899\
        );

    \I__14976\ : InMux
    port map (
            O => \N__60978\,
            I => \N__60894\
        );

    \I__14975\ : InMux
    port map (
            O => \N__60977\,
            I => \N__60894\
        );

    \I__14974\ : InMux
    port map (
            O => \N__60976\,
            I => \N__60889\
        );

    \I__14973\ : InMux
    port map (
            O => \N__60975\,
            I => \N__60889\
        );

    \I__14972\ : LocalMux
    port map (
            O => \N__60970\,
            I => \N__60884\
        );

    \I__14971\ : LocalMux
    port map (
            O => \N__60963\,
            I => \N__60884\
        );

    \I__14970\ : LocalMux
    port map (
            O => \N__60958\,
            I => \N__60881\
        );

    \I__14969\ : InMux
    port map (
            O => \N__60957\,
            I => \N__60876\
        );

    \I__14968\ : InMux
    port map (
            O => \N__60956\,
            I => \N__60871\
        );

    \I__14967\ : InMux
    port map (
            O => \N__60955\,
            I => \N__60871\
        );

    \I__14966\ : InMux
    port map (
            O => \N__60954\,
            I => \N__60866\
        );

    \I__14965\ : InMux
    port map (
            O => \N__60953\,
            I => \N__60866\
        );

    \I__14964\ : InMux
    port map (
            O => \N__60952\,
            I => \N__60862\
        );

    \I__14963\ : InMux
    port map (
            O => \N__60949\,
            I => \N__60859\
        );

    \I__14962\ : InMux
    port map (
            O => \N__60948\,
            I => \N__60856\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__60945\,
            I => \N__60853\
        );

    \I__14960\ : Span12Mux_v
    port map (
            O => \N__60942\,
            I => \N__60850\
        );

    \I__14959\ : LocalMux
    port map (
            O => \N__60939\,
            I => \N__60847\
        );

    \I__14958\ : Span4Mux_h
    port map (
            O => \N__60932\,
            I => \N__60842\
        );

    \I__14957\ : Span4Mux_h
    port map (
            O => \N__60929\,
            I => \N__60842\
        );

    \I__14956\ : LocalMux
    port map (
            O => \N__60926\,
            I => \N__60837\
        );

    \I__14955\ : LocalMux
    port map (
            O => \N__60921\,
            I => \N__60837\
        );

    \I__14954\ : LocalMux
    port map (
            O => \N__60918\,
            I => \N__60834\
        );

    \I__14953\ : LocalMux
    port map (
            O => \N__60915\,
            I => \N__60831\
        );

    \I__14952\ : LocalMux
    port map (
            O => \N__60912\,
            I => \N__60822\
        );

    \I__14951\ : Span4Mux_v
    port map (
            O => \N__60909\,
            I => \N__60822\
        );

    \I__14950\ : Span4Mux_h
    port map (
            O => \N__60906\,
            I => \N__60822\
        );

    \I__14949\ : LocalMux
    port map (
            O => \N__60903\,
            I => \N__60822\
        );

    \I__14948\ : InMux
    port map (
            O => \N__60902\,
            I => \N__60819\
        );

    \I__14947\ : LocalMux
    port map (
            O => \N__60899\,
            I => \N__60810\
        );

    \I__14946\ : LocalMux
    port map (
            O => \N__60894\,
            I => \N__60810\
        );

    \I__14945\ : LocalMux
    port map (
            O => \N__60889\,
            I => \N__60810\
        );

    \I__14944\ : Span4Mux_v
    port map (
            O => \N__60884\,
            I => \N__60810\
        );

    \I__14943\ : Span4Mux_h
    port map (
            O => \N__60881\,
            I => \N__60807\
        );

    \I__14942\ : InMux
    port map (
            O => \N__60880\,
            I => \N__60804\
        );

    \I__14941\ : InMux
    port map (
            O => \N__60879\,
            I => \N__60801\
        );

    \I__14940\ : LocalMux
    port map (
            O => \N__60876\,
            I => \N__60794\
        );

    \I__14939\ : LocalMux
    port map (
            O => \N__60871\,
            I => \N__60794\
        );

    \I__14938\ : LocalMux
    port map (
            O => \N__60866\,
            I => \N__60794\
        );

    \I__14937\ : InMux
    port map (
            O => \N__60865\,
            I => \N__60789\
        );

    \I__14936\ : LocalMux
    port map (
            O => \N__60862\,
            I => \N__60786\
        );

    \I__14935\ : LocalMux
    port map (
            O => \N__60859\,
            I => \N__60781\
        );

    \I__14934\ : LocalMux
    port map (
            O => \N__60856\,
            I => \N__60781\
        );

    \I__14933\ : Span12Mux_h
    port map (
            O => \N__60853\,
            I => \N__60778\
        );

    \I__14932\ : Span12Mux_h
    port map (
            O => \N__60850\,
            I => \N__60775\
        );

    \I__14931\ : Span4Mux_h
    port map (
            O => \N__60847\,
            I => \N__60770\
        );

    \I__14930\ : Span4Mux_h
    port map (
            O => \N__60842\,
            I => \N__60770\
        );

    \I__14929\ : Span4Mux_v
    port map (
            O => \N__60837\,
            I => \N__60757\
        );

    \I__14928\ : Span4Mux_v
    port map (
            O => \N__60834\,
            I => \N__60757\
        );

    \I__14927\ : Span4Mux_v
    port map (
            O => \N__60831\,
            I => \N__60757\
        );

    \I__14926\ : Span4Mux_h
    port map (
            O => \N__60822\,
            I => \N__60757\
        );

    \I__14925\ : LocalMux
    port map (
            O => \N__60819\,
            I => \N__60757\
        );

    \I__14924\ : Span4Mux_v
    port map (
            O => \N__60810\,
            I => \N__60757\
        );

    \I__14923\ : Span4Mux_h
    port map (
            O => \N__60807\,
            I => \N__60750\
        );

    \I__14922\ : LocalMux
    port map (
            O => \N__60804\,
            I => \N__60750\
        );

    \I__14921\ : LocalMux
    port map (
            O => \N__60801\,
            I => \N__60750\
        );

    \I__14920\ : Span4Mux_v
    port map (
            O => \N__60794\,
            I => \N__60747\
        );

    \I__14919\ : InMux
    port map (
            O => \N__60793\,
            I => \N__60742\
        );

    \I__14918\ : InMux
    port map (
            O => \N__60792\,
            I => \N__60742\
        );

    \I__14917\ : LocalMux
    port map (
            O => \N__60789\,
            I => comm_cmd_3
        );

    \I__14916\ : Odrv4
    port map (
            O => \N__60786\,
            I => comm_cmd_3
        );

    \I__14915\ : Odrv12
    port map (
            O => \N__60781\,
            I => comm_cmd_3
        );

    \I__14914\ : Odrv12
    port map (
            O => \N__60778\,
            I => comm_cmd_3
        );

    \I__14913\ : Odrv12
    port map (
            O => \N__60775\,
            I => comm_cmd_3
        );

    \I__14912\ : Odrv4
    port map (
            O => \N__60770\,
            I => comm_cmd_3
        );

    \I__14911\ : Odrv4
    port map (
            O => \N__60757\,
            I => comm_cmd_3
        );

    \I__14910\ : Odrv4
    port map (
            O => \N__60750\,
            I => comm_cmd_3
        );

    \I__14909\ : Odrv4
    port map (
            O => \N__60747\,
            I => comm_cmd_3
        );

    \I__14908\ : LocalMux
    port map (
            O => \N__60742\,
            I => comm_cmd_3
        );

    \I__14907\ : InMux
    port map (
            O => \N__60721\,
            I => \N__60718\
        );

    \I__14906\ : LocalMux
    port map (
            O => \N__60718\,
            I => \N__60715\
        );

    \I__14905\ : Odrv4
    port map (
            O => \N__60715\,
            I => n23492
        );

    \I__14904\ : CascadeMux
    port map (
            O => \N__60712\,
            I => \N__60709\
        );

    \I__14903\ : InMux
    port map (
            O => \N__60709\,
            I => \N__60706\
        );

    \I__14902\ : LocalMux
    port map (
            O => \N__60706\,
            I => \N__60703\
        );

    \I__14901\ : Sp12to4
    port map (
            O => \N__60703\,
            I => \N__60700\
        );

    \I__14900\ : Odrv12
    port map (
            O => \N__60700\,
            I => n23_adj_1773
        );

    \I__14899\ : InMux
    port map (
            O => \N__60697\,
            I => \N__60694\
        );

    \I__14898\ : LocalMux
    port map (
            O => \N__60694\,
            I => \N__60691\
        );

    \I__14897\ : Span12Mux_h
    port map (
            O => \N__60691\,
            I => \N__60686\
        );

    \I__14896\ : InMux
    port map (
            O => \N__60690\,
            I => \N__60681\
        );

    \I__14895\ : InMux
    port map (
            O => \N__60689\,
            I => \N__60681\
        );

    \I__14894\ : Odrv12
    port map (
            O => \N__60686\,
            I => req_data_cnt_13
        );

    \I__14893\ : LocalMux
    port map (
            O => \N__60681\,
            I => req_data_cnt_13
        );

    \I__14892\ : InMux
    port map (
            O => \N__60676\,
            I => \N__60673\
        );

    \I__14891\ : LocalMux
    port map (
            O => \N__60673\,
            I => n25_adj_1774
        );

    \I__14890\ : InMux
    port map (
            O => \N__60670\,
            I => \N__60660\
        );

    \I__14889\ : InMux
    port map (
            O => \N__60669\,
            I => \N__60657\
        );

    \I__14888\ : InMux
    port map (
            O => \N__60668\,
            I => \N__60650\
        );

    \I__14887\ : InMux
    port map (
            O => \N__60667\,
            I => \N__60650\
        );

    \I__14886\ : InMux
    port map (
            O => \N__60666\,
            I => \N__60650\
        );

    \I__14885\ : InMux
    port map (
            O => \N__60665\,
            I => \N__60643\
        );

    \I__14884\ : InMux
    port map (
            O => \N__60664\,
            I => \N__60637\
        );

    \I__14883\ : CascadeMux
    port map (
            O => \N__60663\,
            I => \N__60632\
        );

    \I__14882\ : LocalMux
    port map (
            O => \N__60660\,
            I => \N__60628\
        );

    \I__14881\ : LocalMux
    port map (
            O => \N__60657\,
            I => \N__60624\
        );

    \I__14880\ : LocalMux
    port map (
            O => \N__60650\,
            I => \N__60621\
        );

    \I__14879\ : InMux
    port map (
            O => \N__60649\,
            I => \N__60616\
        );

    \I__14878\ : InMux
    port map (
            O => \N__60648\,
            I => \N__60612\
        );

    \I__14877\ : InMux
    port map (
            O => \N__60647\,
            I => \N__60604\
        );

    \I__14876\ : InMux
    port map (
            O => \N__60646\,
            I => \N__60604\
        );

    \I__14875\ : LocalMux
    port map (
            O => \N__60643\,
            I => \N__60584\
        );

    \I__14874\ : InMux
    port map (
            O => \N__60642\,
            I => \N__60579\
        );

    \I__14873\ : InMux
    port map (
            O => \N__60641\,
            I => \N__60579\
        );

    \I__14872\ : InMux
    port map (
            O => \N__60640\,
            I => \N__60576\
        );

    \I__14871\ : LocalMux
    port map (
            O => \N__60637\,
            I => \N__60573\
        );

    \I__14870\ : InMux
    port map (
            O => \N__60636\,
            I => \N__60568\
        );

    \I__14869\ : InMux
    port map (
            O => \N__60635\,
            I => \N__60568\
        );

    \I__14868\ : InMux
    port map (
            O => \N__60632\,
            I => \N__60565\
        );

    \I__14867\ : InMux
    port map (
            O => \N__60631\,
            I => \N__60561\
        );

    \I__14866\ : Span4Mux_h
    port map (
            O => \N__60628\,
            I => \N__60558\
        );

    \I__14865\ : InMux
    port map (
            O => \N__60627\,
            I => \N__60555\
        );

    \I__14864\ : Span4Mux_h
    port map (
            O => \N__60624\,
            I => \N__60550\
        );

    \I__14863\ : Span4Mux_h
    port map (
            O => \N__60621\,
            I => \N__60550\
        );

    \I__14862\ : InMux
    port map (
            O => \N__60620\,
            I => \N__60547\
        );

    \I__14861\ : InMux
    port map (
            O => \N__60619\,
            I => \N__60540\
        );

    \I__14860\ : LocalMux
    port map (
            O => \N__60616\,
            I => \N__60537\
        );

    \I__14859\ : InMux
    port map (
            O => \N__60615\,
            I => \N__60534\
        );

    \I__14858\ : LocalMux
    port map (
            O => \N__60612\,
            I => \N__60531\
        );

    \I__14857\ : InMux
    port map (
            O => \N__60611\,
            I => \N__60528\
        );

    \I__14856\ : InMux
    port map (
            O => \N__60610\,
            I => \N__60523\
        );

    \I__14855\ : InMux
    port map (
            O => \N__60609\,
            I => \N__60523\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__60604\,
            I => \N__60513\
        );

    \I__14853\ : InMux
    port map (
            O => \N__60603\,
            I => \N__60510\
        );

    \I__14852\ : InMux
    port map (
            O => \N__60602\,
            I => \N__60507\
        );

    \I__14851\ : InMux
    port map (
            O => \N__60601\,
            I => \N__60502\
        );

    \I__14850\ : InMux
    port map (
            O => \N__60600\,
            I => \N__60502\
        );

    \I__14849\ : InMux
    port map (
            O => \N__60599\,
            I => \N__60490\
        );

    \I__14848\ : InMux
    port map (
            O => \N__60598\,
            I => \N__60490\
        );

    \I__14847\ : InMux
    port map (
            O => \N__60597\,
            I => \N__60487\
        );

    \I__14846\ : InMux
    port map (
            O => \N__60596\,
            I => \N__60480\
        );

    \I__14845\ : InMux
    port map (
            O => \N__60595\,
            I => \N__60480\
        );

    \I__14844\ : InMux
    port map (
            O => \N__60594\,
            I => \N__60480\
        );

    \I__14843\ : InMux
    port map (
            O => \N__60593\,
            I => \N__60475\
        );

    \I__14842\ : InMux
    port map (
            O => \N__60592\,
            I => \N__60470\
        );

    \I__14841\ : InMux
    port map (
            O => \N__60591\,
            I => \N__60470\
        );

    \I__14840\ : InMux
    port map (
            O => \N__60590\,
            I => \N__60464\
        );

    \I__14839\ : InMux
    port map (
            O => \N__60589\,
            I => \N__60458\
        );

    \I__14838\ : InMux
    port map (
            O => \N__60588\,
            I => \N__60453\
        );

    \I__14837\ : InMux
    port map (
            O => \N__60587\,
            I => \N__60453\
        );

    \I__14836\ : Span4Mux_h
    port map (
            O => \N__60584\,
            I => \N__60446\
        );

    \I__14835\ : LocalMux
    port map (
            O => \N__60579\,
            I => \N__60446\
        );

    \I__14834\ : LocalMux
    port map (
            O => \N__60576\,
            I => \N__60446\
        );

    \I__14833\ : Span4Mux_v
    port map (
            O => \N__60573\,
            I => \N__60439\
        );

    \I__14832\ : LocalMux
    port map (
            O => \N__60568\,
            I => \N__60439\
        );

    \I__14831\ : LocalMux
    port map (
            O => \N__60565\,
            I => \N__60439\
        );

    \I__14830\ : InMux
    port map (
            O => \N__60564\,
            I => \N__60436\
        );

    \I__14829\ : LocalMux
    port map (
            O => \N__60561\,
            I => \N__60433\
        );

    \I__14828\ : Span4Mux_h
    port map (
            O => \N__60558\,
            I => \N__60426\
        );

    \I__14827\ : LocalMux
    port map (
            O => \N__60555\,
            I => \N__60426\
        );

    \I__14826\ : Span4Mux_h
    port map (
            O => \N__60550\,
            I => \N__60426\
        );

    \I__14825\ : LocalMux
    port map (
            O => \N__60547\,
            I => \N__60423\
        );

    \I__14824\ : InMux
    port map (
            O => \N__60546\,
            I => \N__60416\
        );

    \I__14823\ : InMux
    port map (
            O => \N__60545\,
            I => \N__60416\
        );

    \I__14822\ : InMux
    port map (
            O => \N__60544\,
            I => \N__60416\
        );

    \I__14821\ : InMux
    port map (
            O => \N__60543\,
            I => \N__60413\
        );

    \I__14820\ : LocalMux
    port map (
            O => \N__60540\,
            I => \N__60410\
        );

    \I__14819\ : Span4Mux_v
    port map (
            O => \N__60537\,
            I => \N__60407\
        );

    \I__14818\ : LocalMux
    port map (
            O => \N__60534\,
            I => \N__60398\
        );

    \I__14817\ : Span4Mux_v
    port map (
            O => \N__60531\,
            I => \N__60398\
        );

    \I__14816\ : LocalMux
    port map (
            O => \N__60528\,
            I => \N__60398\
        );

    \I__14815\ : LocalMux
    port map (
            O => \N__60523\,
            I => \N__60398\
        );

    \I__14814\ : InMux
    port map (
            O => \N__60522\,
            I => \N__60392\
        );

    \I__14813\ : InMux
    port map (
            O => \N__60521\,
            I => \N__60389\
        );

    \I__14812\ : InMux
    port map (
            O => \N__60520\,
            I => \N__60386\
        );

    \I__14811\ : InMux
    port map (
            O => \N__60519\,
            I => \N__60381\
        );

    \I__14810\ : InMux
    port map (
            O => \N__60518\,
            I => \N__60381\
        );

    \I__14809\ : InMux
    port map (
            O => \N__60517\,
            I => \N__60376\
        );

    \I__14808\ : InMux
    port map (
            O => \N__60516\,
            I => \N__60376\
        );

    \I__14807\ : Span4Mux_h
    port map (
            O => \N__60513\,
            I => \N__60371\
        );

    \I__14806\ : LocalMux
    port map (
            O => \N__60510\,
            I => \N__60371\
        );

    \I__14805\ : LocalMux
    port map (
            O => \N__60507\,
            I => \N__60366\
        );

    \I__14804\ : LocalMux
    port map (
            O => \N__60502\,
            I => \N__60366\
        );

    \I__14803\ : InMux
    port map (
            O => \N__60501\,
            I => \N__60359\
        );

    \I__14802\ : InMux
    port map (
            O => \N__60500\,
            I => \N__60359\
        );

    \I__14801\ : InMux
    port map (
            O => \N__60499\,
            I => \N__60359\
        );

    \I__14800\ : InMux
    port map (
            O => \N__60498\,
            I => \N__60354\
        );

    \I__14799\ : InMux
    port map (
            O => \N__60497\,
            I => \N__60349\
        );

    \I__14798\ : InMux
    port map (
            O => \N__60496\,
            I => \N__60344\
        );

    \I__14797\ : InMux
    port map (
            O => \N__60495\,
            I => \N__60344\
        );

    \I__14796\ : LocalMux
    port map (
            O => \N__60490\,
            I => \N__60341\
        );

    \I__14795\ : LocalMux
    port map (
            O => \N__60487\,
            I => \N__60336\
        );

    \I__14794\ : LocalMux
    port map (
            O => \N__60480\,
            I => \N__60336\
        );

    \I__14793\ : InMux
    port map (
            O => \N__60479\,
            I => \N__60331\
        );

    \I__14792\ : InMux
    port map (
            O => \N__60478\,
            I => \N__60331\
        );

    \I__14791\ : LocalMux
    port map (
            O => \N__60475\,
            I => \N__60326\
        );

    \I__14790\ : LocalMux
    port map (
            O => \N__60470\,
            I => \N__60326\
        );

    \I__14789\ : InMux
    port map (
            O => \N__60469\,
            I => \N__60321\
        );

    \I__14788\ : InMux
    port map (
            O => \N__60468\,
            I => \N__60321\
        );

    \I__14787\ : InMux
    port map (
            O => \N__60467\,
            I => \N__60318\
        );

    \I__14786\ : LocalMux
    port map (
            O => \N__60464\,
            I => \N__60315\
        );

    \I__14785\ : CascadeMux
    port map (
            O => \N__60463\,
            I => \N__60310\
        );

    \I__14784\ : InMux
    port map (
            O => \N__60462\,
            I => \N__60304\
        );

    \I__14783\ : InMux
    port map (
            O => \N__60461\,
            I => \N__60304\
        );

    \I__14782\ : LocalMux
    port map (
            O => \N__60458\,
            I => \N__60301\
        );

    \I__14781\ : LocalMux
    port map (
            O => \N__60453\,
            I => \N__60294\
        );

    \I__14780\ : Span4Mux_h
    port map (
            O => \N__60446\,
            I => \N__60294\
        );

    \I__14779\ : Span4Mux_h
    port map (
            O => \N__60439\,
            I => \N__60294\
        );

    \I__14778\ : LocalMux
    port map (
            O => \N__60436\,
            I => \N__60285\
        );

    \I__14777\ : Span4Mux_h
    port map (
            O => \N__60433\,
            I => \N__60285\
        );

    \I__14776\ : Span4Mux_v
    port map (
            O => \N__60426\,
            I => \N__60285\
        );

    \I__14775\ : Span4Mux_h
    port map (
            O => \N__60423\,
            I => \N__60285\
        );

    \I__14774\ : LocalMux
    port map (
            O => \N__60416\,
            I => \N__60282\
        );

    \I__14773\ : LocalMux
    port map (
            O => \N__60413\,
            I => \N__60273\
        );

    \I__14772\ : Span4Mux_h
    port map (
            O => \N__60410\,
            I => \N__60273\
        );

    \I__14771\ : Span4Mux_v
    port map (
            O => \N__60407\,
            I => \N__60273\
        );

    \I__14770\ : Span4Mux_v
    port map (
            O => \N__60398\,
            I => \N__60273\
        );

    \I__14769\ : CascadeMux
    port map (
            O => \N__60397\,
            I => \N__60270\
        );

    \I__14768\ : InMux
    port map (
            O => \N__60396\,
            I => \N__60266\
        );

    \I__14767\ : InMux
    port map (
            O => \N__60395\,
            I => \N__60263\
        );

    \I__14766\ : LocalMux
    port map (
            O => \N__60392\,
            I => \N__60251\
        );

    \I__14765\ : LocalMux
    port map (
            O => \N__60389\,
            I => \N__60251\
        );

    \I__14764\ : LocalMux
    port map (
            O => \N__60386\,
            I => \N__60251\
        );

    \I__14763\ : LocalMux
    port map (
            O => \N__60381\,
            I => \N__60251\
        );

    \I__14762\ : LocalMux
    port map (
            O => \N__60376\,
            I => \N__60251\
        );

    \I__14761\ : Span4Mux_v
    port map (
            O => \N__60371\,
            I => \N__60240\
        );

    \I__14760\ : Span4Mux_v
    port map (
            O => \N__60366\,
            I => \N__60240\
        );

    \I__14759\ : LocalMux
    port map (
            O => \N__60359\,
            I => \N__60240\
        );

    \I__14758\ : InMux
    port map (
            O => \N__60358\,
            I => \N__60237\
        );

    \I__14757\ : CascadeMux
    port map (
            O => \N__60357\,
            I => \N__60234\
        );

    \I__14756\ : LocalMux
    port map (
            O => \N__60354\,
            I => \N__60230\
        );

    \I__14755\ : InMux
    port map (
            O => \N__60353\,
            I => \N__60225\
        );

    \I__14754\ : InMux
    port map (
            O => \N__60352\,
            I => \N__60225\
        );

    \I__14753\ : LocalMux
    port map (
            O => \N__60349\,
            I => \N__60212\
        );

    \I__14752\ : LocalMux
    port map (
            O => \N__60344\,
            I => \N__60212\
        );

    \I__14751\ : Span4Mux_h
    port map (
            O => \N__60341\,
            I => \N__60212\
        );

    \I__14750\ : Span4Mux_h
    port map (
            O => \N__60336\,
            I => \N__60212\
        );

    \I__14749\ : LocalMux
    port map (
            O => \N__60331\,
            I => \N__60212\
        );

    \I__14748\ : Span4Mux_h
    port map (
            O => \N__60326\,
            I => \N__60212\
        );

    \I__14747\ : LocalMux
    port map (
            O => \N__60321\,
            I => \N__60209\
        );

    \I__14746\ : LocalMux
    port map (
            O => \N__60318\,
            I => \N__60204\
        );

    \I__14745\ : Span4Mux_v
    port map (
            O => \N__60315\,
            I => \N__60204\
        );

    \I__14744\ : InMux
    port map (
            O => \N__60314\,
            I => \N__60195\
        );

    \I__14743\ : InMux
    port map (
            O => \N__60313\,
            I => \N__60195\
        );

    \I__14742\ : InMux
    port map (
            O => \N__60310\,
            I => \N__60195\
        );

    \I__14741\ : InMux
    port map (
            O => \N__60309\,
            I => \N__60195\
        );

    \I__14740\ : LocalMux
    port map (
            O => \N__60304\,
            I => \N__60186\
        );

    \I__14739\ : Sp12to4
    port map (
            O => \N__60301\,
            I => \N__60186\
        );

    \I__14738\ : Sp12to4
    port map (
            O => \N__60294\,
            I => \N__60186\
        );

    \I__14737\ : Sp12to4
    port map (
            O => \N__60285\,
            I => \N__60186\
        );

    \I__14736\ : Span4Mux_v
    port map (
            O => \N__60282\,
            I => \N__60181\
        );

    \I__14735\ : Span4Mux_h
    port map (
            O => \N__60273\,
            I => \N__60181\
        );

    \I__14734\ : InMux
    port map (
            O => \N__60270\,
            I => \N__60176\
        );

    \I__14733\ : InMux
    port map (
            O => \N__60269\,
            I => \N__60176\
        );

    \I__14732\ : LocalMux
    port map (
            O => \N__60266\,
            I => \N__60173\
        );

    \I__14731\ : LocalMux
    port map (
            O => \N__60263\,
            I => \N__60170\
        );

    \I__14730\ : InMux
    port map (
            O => \N__60262\,
            I => \N__60167\
        );

    \I__14729\ : Span4Mux_v
    port map (
            O => \N__60251\,
            I => \N__60164\
        );

    \I__14728\ : InMux
    port map (
            O => \N__60250\,
            I => \N__60157\
        );

    \I__14727\ : InMux
    port map (
            O => \N__60249\,
            I => \N__60157\
        );

    \I__14726\ : InMux
    port map (
            O => \N__60248\,
            I => \N__60157\
        );

    \I__14725\ : InMux
    port map (
            O => \N__60247\,
            I => \N__60154\
        );

    \I__14724\ : Span4Mux_h
    port map (
            O => \N__60240\,
            I => \N__60151\
        );

    \I__14723\ : LocalMux
    port map (
            O => \N__60237\,
            I => \N__60148\
        );

    \I__14722\ : InMux
    port map (
            O => \N__60234\,
            I => \N__60143\
        );

    \I__14721\ : InMux
    port map (
            O => \N__60233\,
            I => \N__60143\
        );

    \I__14720\ : Span4Mux_v
    port map (
            O => \N__60230\,
            I => \N__60132\
        );

    \I__14719\ : LocalMux
    port map (
            O => \N__60225\,
            I => \N__60132\
        );

    \I__14718\ : Span4Mux_v
    port map (
            O => \N__60212\,
            I => \N__60132\
        );

    \I__14717\ : Span4Mux_h
    port map (
            O => \N__60209\,
            I => \N__60132\
        );

    \I__14716\ : Span4Mux_h
    port map (
            O => \N__60204\,
            I => \N__60132\
        );

    \I__14715\ : LocalMux
    port map (
            O => \N__60195\,
            I => \N__60123\
        );

    \I__14714\ : Span12Mux_v
    port map (
            O => \N__60186\,
            I => \N__60123\
        );

    \I__14713\ : Sp12to4
    port map (
            O => \N__60181\,
            I => \N__60123\
        );

    \I__14712\ : LocalMux
    port map (
            O => \N__60176\,
            I => \N__60123\
        );

    \I__14711\ : Odrv4
    port map (
            O => \N__60173\,
            I => comm_cmd_1
        );

    \I__14710\ : Odrv12
    port map (
            O => \N__60170\,
            I => comm_cmd_1
        );

    \I__14709\ : LocalMux
    port map (
            O => \N__60167\,
            I => comm_cmd_1
        );

    \I__14708\ : Odrv4
    port map (
            O => \N__60164\,
            I => comm_cmd_1
        );

    \I__14707\ : LocalMux
    port map (
            O => \N__60157\,
            I => comm_cmd_1
        );

    \I__14706\ : LocalMux
    port map (
            O => \N__60154\,
            I => comm_cmd_1
        );

    \I__14705\ : Odrv4
    port map (
            O => \N__60151\,
            I => comm_cmd_1
        );

    \I__14704\ : Odrv12
    port map (
            O => \N__60148\,
            I => comm_cmd_1
        );

    \I__14703\ : LocalMux
    port map (
            O => \N__60143\,
            I => comm_cmd_1
        );

    \I__14702\ : Odrv4
    port map (
            O => \N__60132\,
            I => comm_cmd_1
        );

    \I__14701\ : Odrv12
    port map (
            O => \N__60123\,
            I => comm_cmd_1
        );

    \I__14700\ : InMux
    port map (
            O => \N__60100\,
            I => \N__60087\
        );

    \I__14699\ : InMux
    port map (
            O => \N__60099\,
            I => \N__60084\
        );

    \I__14698\ : InMux
    port map (
            O => \N__60098\,
            I => \N__60077\
        );

    \I__14697\ : CascadeMux
    port map (
            O => \N__60097\,
            I => \N__60073\
        );

    \I__14696\ : InMux
    port map (
            O => \N__60096\,
            I => \N__60069\
        );

    \I__14695\ : InMux
    port map (
            O => \N__60095\,
            I => \N__60066\
        );

    \I__14694\ : InMux
    port map (
            O => \N__60094\,
            I => \N__60060\
        );

    \I__14693\ : InMux
    port map (
            O => \N__60093\,
            I => \N__60053\
        );

    \I__14692\ : InMux
    port map (
            O => \N__60092\,
            I => \N__60053\
        );

    \I__14691\ : CascadeMux
    port map (
            O => \N__60091\,
            I => \N__60049\
        );

    \I__14690\ : CascadeMux
    port map (
            O => \N__60090\,
            I => \N__60037\
        );

    \I__14689\ : LocalMux
    port map (
            O => \N__60087\,
            I => \N__60031\
        );

    \I__14688\ : LocalMux
    port map (
            O => \N__60084\,
            I => \N__60031\
        );

    \I__14687\ : InMux
    port map (
            O => \N__60083\,
            I => \N__60026\
        );

    \I__14686\ : InMux
    port map (
            O => \N__60082\,
            I => \N__60026\
        );

    \I__14685\ : InMux
    port map (
            O => \N__60081\,
            I => \N__60021\
        );

    \I__14684\ : InMux
    port map (
            O => \N__60080\,
            I => \N__60021\
        );

    \I__14683\ : LocalMux
    port map (
            O => \N__60077\,
            I => \N__60018\
        );

    \I__14682\ : InMux
    port map (
            O => \N__60076\,
            I => \N__60015\
        );

    \I__14681\ : InMux
    port map (
            O => \N__60073\,
            I => \N__60009\
        );

    \I__14680\ : InMux
    port map (
            O => \N__60072\,
            I => \N__60009\
        );

    \I__14679\ : LocalMux
    port map (
            O => \N__60069\,
            I => \N__60003\
        );

    \I__14678\ : LocalMux
    port map (
            O => \N__60066\,
            I => \N__59996\
        );

    \I__14677\ : InMux
    port map (
            O => \N__60065\,
            I => \N__59988\
        );

    \I__14676\ : InMux
    port map (
            O => \N__60064\,
            I => \N__59979\
        );

    \I__14675\ : InMux
    port map (
            O => \N__60063\,
            I => \N__59970\
        );

    \I__14674\ : LocalMux
    port map (
            O => \N__60060\,
            I => \N__59966\
        );

    \I__14673\ : InMux
    port map (
            O => \N__60059\,
            I => \N__59955\
        );

    \I__14672\ : InMux
    port map (
            O => \N__60058\,
            I => \N__59955\
        );

    \I__14671\ : LocalMux
    port map (
            O => \N__60053\,
            I => \N__59951\
        );

    \I__14670\ : InMux
    port map (
            O => \N__60052\,
            I => \N__59944\
        );

    \I__14669\ : InMux
    port map (
            O => \N__60049\,
            I => \N__59944\
        );

    \I__14668\ : InMux
    port map (
            O => \N__60048\,
            I => \N__59944\
        );

    \I__14667\ : InMux
    port map (
            O => \N__60047\,
            I => \N__59937\
        );

    \I__14666\ : InMux
    port map (
            O => \N__60046\,
            I => \N__59937\
        );

    \I__14665\ : InMux
    port map (
            O => \N__60045\,
            I => \N__59937\
        );

    \I__14664\ : CascadeMux
    port map (
            O => \N__60044\,
            I => \N__59933\
        );

    \I__14663\ : CascadeMux
    port map (
            O => \N__60043\,
            I => \N__59930\
        );

    \I__14662\ : InMux
    port map (
            O => \N__60042\,
            I => \N__59925\
        );

    \I__14661\ : InMux
    port map (
            O => \N__60041\,
            I => \N__59925\
        );

    \I__14660\ : InMux
    port map (
            O => \N__60040\,
            I => \N__59922\
        );

    \I__14659\ : InMux
    port map (
            O => \N__60037\,
            I => \N__59917\
        );

    \I__14658\ : InMux
    port map (
            O => \N__60036\,
            I => \N__59917\
        );

    \I__14657\ : Span4Mux_v
    port map (
            O => \N__60031\,
            I => \N__59912\
        );

    \I__14656\ : LocalMux
    port map (
            O => \N__60026\,
            I => \N__59912\
        );

    \I__14655\ : LocalMux
    port map (
            O => \N__60021\,
            I => \N__59905\
        );

    \I__14654\ : Span4Mux_v
    port map (
            O => \N__60018\,
            I => \N__59905\
        );

    \I__14653\ : LocalMux
    port map (
            O => \N__60015\,
            I => \N__59905\
        );

    \I__14652\ : CascadeMux
    port map (
            O => \N__60014\,
            I => \N__59901\
        );

    \I__14651\ : LocalMux
    port map (
            O => \N__60009\,
            I => \N__59897\
        );

    \I__14650\ : InMux
    port map (
            O => \N__60008\,
            I => \N__59894\
        );

    \I__14649\ : InMux
    port map (
            O => \N__60007\,
            I => \N__59891\
        );

    \I__14648\ : InMux
    port map (
            O => \N__60006\,
            I => \N__59888\
        );

    \I__14647\ : Span4Mux_v
    port map (
            O => \N__60003\,
            I => \N__59884\
        );

    \I__14646\ : InMux
    port map (
            O => \N__60002\,
            I => \N__59881\
        );

    \I__14645\ : InMux
    port map (
            O => \N__60001\,
            I => \N__59874\
        );

    \I__14644\ : InMux
    port map (
            O => \N__60000\,
            I => \N__59874\
        );

    \I__14643\ : InMux
    port map (
            O => \N__59999\,
            I => \N__59874\
        );

    \I__14642\ : Span4Mux_v
    port map (
            O => \N__59996\,
            I => \N__59871\
        );

    \I__14641\ : InMux
    port map (
            O => \N__59995\,
            I => \N__59868\
        );

    \I__14640\ : InMux
    port map (
            O => \N__59994\,
            I => \N__59862\
        );

    \I__14639\ : InMux
    port map (
            O => \N__59993\,
            I => \N__59862\
        );

    \I__14638\ : InMux
    port map (
            O => \N__59992\,
            I => \N__59857\
        );

    \I__14637\ : InMux
    port map (
            O => \N__59991\,
            I => \N__59857\
        );

    \I__14636\ : LocalMux
    port map (
            O => \N__59988\,
            I => \N__59854\
        );

    \I__14635\ : InMux
    port map (
            O => \N__59987\,
            I => \N__59851\
        );

    \I__14634\ : InMux
    port map (
            O => \N__59986\,
            I => \N__59846\
        );

    \I__14633\ : InMux
    port map (
            O => \N__59985\,
            I => \N__59846\
        );

    \I__14632\ : InMux
    port map (
            O => \N__59984\,
            I => \N__59839\
        );

    \I__14631\ : InMux
    port map (
            O => \N__59983\,
            I => \N__59839\
        );

    \I__14630\ : InMux
    port map (
            O => \N__59982\,
            I => \N__59839\
        );

    \I__14629\ : LocalMux
    port map (
            O => \N__59979\,
            I => \N__59836\
        );

    \I__14628\ : InMux
    port map (
            O => \N__59978\,
            I => \N__59831\
        );

    \I__14627\ : InMux
    port map (
            O => \N__59977\,
            I => \N__59831\
        );

    \I__14626\ : InMux
    port map (
            O => \N__59976\,
            I => \N__59828\
        );

    \I__14625\ : InMux
    port map (
            O => \N__59975\,
            I => \N__59823\
        );

    \I__14624\ : InMux
    port map (
            O => \N__59974\,
            I => \N__59823\
        );

    \I__14623\ : CascadeMux
    port map (
            O => \N__59973\,
            I => \N__59819\
        );

    \I__14622\ : LocalMux
    port map (
            O => \N__59970\,
            I => \N__59816\
        );

    \I__14621\ : InMux
    port map (
            O => \N__59969\,
            I => \N__59813\
        );

    \I__14620\ : Span4Mux_h
    port map (
            O => \N__59966\,
            I => \N__59809\
        );

    \I__14619\ : InMux
    port map (
            O => \N__59965\,
            I => \N__59802\
        );

    \I__14618\ : InMux
    port map (
            O => \N__59964\,
            I => \N__59802\
        );

    \I__14617\ : InMux
    port map (
            O => \N__59963\,
            I => \N__59802\
        );

    \I__14616\ : InMux
    port map (
            O => \N__59962\,
            I => \N__59797\
        );

    \I__14615\ : InMux
    port map (
            O => \N__59961\,
            I => \N__59797\
        );

    \I__14614\ : InMux
    port map (
            O => \N__59960\,
            I => \N__59794\
        );

    \I__14613\ : LocalMux
    port map (
            O => \N__59955\,
            I => \N__59791\
        );

    \I__14612\ : InMux
    port map (
            O => \N__59954\,
            I => \N__59788\
        );

    \I__14611\ : Span4Mux_v
    port map (
            O => \N__59951\,
            I => \N__59785\
        );

    \I__14610\ : LocalMux
    port map (
            O => \N__59944\,
            I => \N__59780\
        );

    \I__14609\ : LocalMux
    port map (
            O => \N__59937\,
            I => \N__59780\
        );

    \I__14608\ : InMux
    port map (
            O => \N__59936\,
            I => \N__59777\
        );

    \I__14607\ : InMux
    port map (
            O => \N__59933\,
            I => \N__59772\
        );

    \I__14606\ : InMux
    port map (
            O => \N__59930\,
            I => \N__59772\
        );

    \I__14605\ : LocalMux
    port map (
            O => \N__59925\,
            I => \N__59769\
        );

    \I__14604\ : LocalMux
    port map (
            O => \N__59922\,
            I => \N__59764\
        );

    \I__14603\ : LocalMux
    port map (
            O => \N__59917\,
            I => \N__59764\
        );

    \I__14602\ : Span4Mux_h
    port map (
            O => \N__59912\,
            I => \N__59759\
        );

    \I__14601\ : Span4Mux_v
    port map (
            O => \N__59905\,
            I => \N__59759\
        );

    \I__14600\ : InMux
    port map (
            O => \N__59904\,
            I => \N__59756\
        );

    \I__14599\ : InMux
    port map (
            O => \N__59901\,
            I => \N__59751\
        );

    \I__14598\ : InMux
    port map (
            O => \N__59900\,
            I => \N__59751\
        );

    \I__14597\ : Span4Mux_h
    port map (
            O => \N__59897\,
            I => \N__59748\
        );

    \I__14596\ : LocalMux
    port map (
            O => \N__59894\,
            I => \N__59743\
        );

    \I__14595\ : LocalMux
    port map (
            O => \N__59891\,
            I => \N__59743\
        );

    \I__14594\ : LocalMux
    port map (
            O => \N__59888\,
            I => \N__59740\
        );

    \I__14593\ : InMux
    port map (
            O => \N__59887\,
            I => \N__59737\
        );

    \I__14592\ : Span4Mux_h
    port map (
            O => \N__59884\,
            I => \N__59734\
        );

    \I__14591\ : LocalMux
    port map (
            O => \N__59881\,
            I => \N__59725\
        );

    \I__14590\ : LocalMux
    port map (
            O => \N__59874\,
            I => \N__59725\
        );

    \I__14589\ : Span4Mux_h
    port map (
            O => \N__59871\,
            I => \N__59725\
        );

    \I__14588\ : LocalMux
    port map (
            O => \N__59868\,
            I => \N__59725\
        );

    \I__14587\ : InMux
    port map (
            O => \N__59867\,
            I => \N__59722\
        );

    \I__14586\ : LocalMux
    port map (
            O => \N__59862\,
            I => \N__59717\
        );

    \I__14585\ : LocalMux
    port map (
            O => \N__59857\,
            I => \N__59717\
        );

    \I__14584\ : Span4Mux_v
    port map (
            O => \N__59854\,
            I => \N__59704\
        );

    \I__14583\ : LocalMux
    port map (
            O => \N__59851\,
            I => \N__59704\
        );

    \I__14582\ : LocalMux
    port map (
            O => \N__59846\,
            I => \N__59704\
        );

    \I__14581\ : LocalMux
    port map (
            O => \N__59839\,
            I => \N__59704\
        );

    \I__14580\ : Span4Mux_h
    port map (
            O => \N__59836\,
            I => \N__59704\
        );

    \I__14579\ : LocalMux
    port map (
            O => \N__59831\,
            I => \N__59704\
        );

    \I__14578\ : LocalMux
    port map (
            O => \N__59828\,
            I => \N__59697\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__59823\,
            I => \N__59697\
        );

    \I__14576\ : InMux
    port map (
            O => \N__59822\,
            I => \N__59692\
        );

    \I__14575\ : InMux
    port map (
            O => \N__59819\,
            I => \N__59692\
        );

    \I__14574\ : Span4Mux_h
    port map (
            O => \N__59816\,
            I => \N__59687\
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__59813\,
            I => \N__59687\
        );

    \I__14572\ : InMux
    port map (
            O => \N__59812\,
            I => \N__59684\
        );

    \I__14571\ : Span4Mux_h
    port map (
            O => \N__59809\,
            I => \N__59673\
        );

    \I__14570\ : LocalMux
    port map (
            O => \N__59802\,
            I => \N__59673\
        );

    \I__14569\ : LocalMux
    port map (
            O => \N__59797\,
            I => \N__59673\
        );

    \I__14568\ : LocalMux
    port map (
            O => \N__59794\,
            I => \N__59673\
        );

    \I__14567\ : Span4Mux_h
    port map (
            O => \N__59791\,
            I => \N__59673\
        );

    \I__14566\ : LocalMux
    port map (
            O => \N__59788\,
            I => \N__59661\
        );

    \I__14565\ : Sp12to4
    port map (
            O => \N__59785\,
            I => \N__59661\
        );

    \I__14564\ : Span12Mux_h
    port map (
            O => \N__59780\,
            I => \N__59661\
        );

    \I__14563\ : LocalMux
    port map (
            O => \N__59777\,
            I => \N__59661\
        );

    \I__14562\ : LocalMux
    port map (
            O => \N__59772\,
            I => \N__59661\
        );

    \I__14561\ : Span4Mux_v
    port map (
            O => \N__59769\,
            I => \N__59654\
        );

    \I__14560\ : Span4Mux_v
    port map (
            O => \N__59764\,
            I => \N__59654\
        );

    \I__14559\ : Span4Mux_h
    port map (
            O => \N__59759\,
            I => \N__59654\
        );

    \I__14558\ : LocalMux
    port map (
            O => \N__59756\,
            I => \N__59649\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__59751\,
            I => \N__59649\
        );

    \I__14556\ : Span4Mux_v
    port map (
            O => \N__59748\,
            I => \N__59644\
        );

    \I__14555\ : Span4Mux_h
    port map (
            O => \N__59743\,
            I => \N__59644\
        );

    \I__14554\ : Span4Mux_v
    port map (
            O => \N__59740\,
            I => \N__59629\
        );

    \I__14553\ : LocalMux
    port map (
            O => \N__59737\,
            I => \N__59629\
        );

    \I__14552\ : Span4Mux_h
    port map (
            O => \N__59734\,
            I => \N__59629\
        );

    \I__14551\ : Span4Mux_v
    port map (
            O => \N__59725\,
            I => \N__59629\
        );

    \I__14550\ : LocalMux
    port map (
            O => \N__59722\,
            I => \N__59629\
        );

    \I__14549\ : Span4Mux_v
    port map (
            O => \N__59717\,
            I => \N__59629\
        );

    \I__14548\ : Span4Mux_v
    port map (
            O => \N__59704\,
            I => \N__59629\
        );

    \I__14547\ : InMux
    port map (
            O => \N__59703\,
            I => \N__59624\
        );

    \I__14546\ : InMux
    port map (
            O => \N__59702\,
            I => \N__59624\
        );

    \I__14545\ : Span4Mux_v
    port map (
            O => \N__59697\,
            I => \N__59619\
        );

    \I__14544\ : LocalMux
    port map (
            O => \N__59692\,
            I => \N__59619\
        );

    \I__14543\ : Span4Mux_v
    port map (
            O => \N__59687\,
            I => \N__59612\
        );

    \I__14542\ : LocalMux
    port map (
            O => \N__59684\,
            I => \N__59612\
        );

    \I__14541\ : Span4Mux_v
    port map (
            O => \N__59673\,
            I => \N__59612\
        );

    \I__14540\ : InMux
    port map (
            O => \N__59672\,
            I => \N__59609\
        );

    \I__14539\ : Span12Mux_h
    port map (
            O => \N__59661\,
            I => \N__59606\
        );

    \I__14538\ : Span4Mux_h
    port map (
            O => \N__59654\,
            I => \N__59601\
        );

    \I__14537\ : Span4Mux_v
    port map (
            O => \N__59649\,
            I => \N__59601\
        );

    \I__14536\ : Odrv4
    port map (
            O => \N__59644\,
            I => comm_cmd_2
        );

    \I__14535\ : Odrv4
    port map (
            O => \N__59629\,
            I => comm_cmd_2
        );

    \I__14534\ : LocalMux
    port map (
            O => \N__59624\,
            I => comm_cmd_2
        );

    \I__14533\ : Odrv4
    port map (
            O => \N__59619\,
            I => comm_cmd_2
        );

    \I__14532\ : Odrv4
    port map (
            O => \N__59612\,
            I => comm_cmd_2
        );

    \I__14531\ : LocalMux
    port map (
            O => \N__59609\,
            I => comm_cmd_2
        );

    \I__14530\ : Odrv12
    port map (
            O => \N__59606\,
            I => comm_cmd_2
        );

    \I__14529\ : Odrv4
    port map (
            O => \N__59601\,
            I => comm_cmd_2
        );

    \I__14528\ : CascadeMux
    port map (
            O => \N__59584\,
            I => \N__59581\
        );

    \I__14527\ : InMux
    port map (
            O => \N__59581\,
            I => \N__59578\
        );

    \I__14526\ : LocalMux
    port map (
            O => \N__59578\,
            I => \N__59575\
        );

    \I__14525\ : Odrv4
    port map (
            O => \N__59575\,
            I => n22316
        );

    \I__14524\ : InMux
    port map (
            O => \N__59572\,
            I => \N__59569\
        );

    \I__14523\ : LocalMux
    port map (
            O => \N__59569\,
            I => n26_adj_1792
        );

    \I__14522\ : InMux
    port map (
            O => \N__59566\,
            I => \N__59563\
        );

    \I__14521\ : LocalMux
    port map (
            O => \N__59563\,
            I => n23456
        );

    \I__14520\ : InMux
    port map (
            O => \N__59560\,
            I => \N__59557\
        );

    \I__14519\ : LocalMux
    port map (
            O => \N__59557\,
            I => buf_data_iac_13
        );

    \I__14518\ : InMux
    port map (
            O => \N__59554\,
            I => \N__59551\
        );

    \I__14517\ : LocalMux
    port map (
            O => \N__59551\,
            I => \N__59548\
        );

    \I__14516\ : Span4Mux_h
    port map (
            O => \N__59548\,
            I => \N__59545\
        );

    \I__14515\ : Odrv4
    port map (
            O => \N__59545\,
            I => n22313
        );

    \I__14514\ : InMux
    port map (
            O => \N__59542\,
            I => \N__59539\
        );

    \I__14513\ : LocalMux
    port map (
            O => \N__59539\,
            I => buf_data_iac_11
        );

    \I__14512\ : InMux
    port map (
            O => \N__59536\,
            I => \N__59533\
        );

    \I__14511\ : LocalMux
    port map (
            O => \N__59533\,
            I => \N__59530\
        );

    \I__14510\ : Odrv12
    port map (
            O => \N__59530\,
            I => n22300
        );

    \I__14509\ : InMux
    port map (
            O => \N__59527\,
            I => \N__59524\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__59524\,
            I => \N__59521\
        );

    \I__14507\ : Odrv4
    port map (
            O => \N__59521\,
            I => buf_data_iac_8
        );

    \I__14506\ : CascadeMux
    port map (
            O => \N__59518\,
            I => \N__59510\
        );

    \I__14505\ : CascadeMux
    port map (
            O => \N__59517\,
            I => \N__59498\
        );

    \I__14504\ : InMux
    port map (
            O => \N__59516\,
            I => \N__59493\
        );

    \I__14503\ : InMux
    port map (
            O => \N__59515\,
            I => \N__59485\
        );

    \I__14502\ : CascadeMux
    port map (
            O => \N__59514\,
            I => \N__59480\
        );

    \I__14501\ : CascadeMux
    port map (
            O => \N__59513\,
            I => \N__59476\
        );

    \I__14500\ : InMux
    port map (
            O => \N__59510\,
            I => \N__59472\
        );

    \I__14499\ : InMux
    port map (
            O => \N__59509\,
            I => \N__59469\
        );

    \I__14498\ : InMux
    port map (
            O => \N__59508\,
            I => \N__59461\
        );

    \I__14497\ : InMux
    port map (
            O => \N__59507\,
            I => \N__59461\
        );

    \I__14496\ : InMux
    port map (
            O => \N__59506\,
            I => \N__59458\
        );

    \I__14495\ : InMux
    port map (
            O => \N__59505\,
            I => \N__59455\
        );

    \I__14494\ : InMux
    port map (
            O => \N__59504\,
            I => \N__59450\
        );

    \I__14493\ : InMux
    port map (
            O => \N__59503\,
            I => \N__59450\
        );

    \I__14492\ : InMux
    port map (
            O => \N__59502\,
            I => \N__59447\
        );

    \I__14491\ : InMux
    port map (
            O => \N__59501\,
            I => \N__59417\
        );

    \I__14490\ : InMux
    port map (
            O => \N__59498\,
            I => \N__59414\
        );

    \I__14489\ : InMux
    port map (
            O => \N__59497\,
            I => \N__59411\
        );

    \I__14488\ : InMux
    port map (
            O => \N__59496\,
            I => \N__59402\
        );

    \I__14487\ : LocalMux
    port map (
            O => \N__59493\,
            I => \N__59394\
        );

    \I__14486\ : InMux
    port map (
            O => \N__59492\,
            I => \N__59391\
        );

    \I__14485\ : InMux
    port map (
            O => \N__59491\,
            I => \N__59388\
        );

    \I__14484\ : InMux
    port map (
            O => \N__59490\,
            I => \N__59381\
        );

    \I__14483\ : InMux
    port map (
            O => \N__59489\,
            I => \N__59381\
        );

    \I__14482\ : InMux
    port map (
            O => \N__59488\,
            I => \N__59381\
        );

    \I__14481\ : LocalMux
    port map (
            O => \N__59485\,
            I => \N__59378\
        );

    \I__14480\ : InMux
    port map (
            O => \N__59484\,
            I => \N__59373\
        );

    \I__14479\ : InMux
    port map (
            O => \N__59483\,
            I => \N__59373\
        );

    \I__14478\ : InMux
    port map (
            O => \N__59480\,
            I => \N__59368\
        );

    \I__14477\ : InMux
    port map (
            O => \N__59479\,
            I => \N__59359\
        );

    \I__14476\ : InMux
    port map (
            O => \N__59476\,
            I => \N__59356\
        );

    \I__14475\ : InMux
    port map (
            O => \N__59475\,
            I => \N__59347\
        );

    \I__14474\ : LocalMux
    port map (
            O => \N__59472\,
            I => \N__59342\
        );

    \I__14473\ : LocalMux
    port map (
            O => \N__59469\,
            I => \N__59342\
        );

    \I__14472\ : InMux
    port map (
            O => \N__59468\,
            I => \N__59337\
        );

    \I__14471\ : InMux
    port map (
            O => \N__59467\,
            I => \N__59337\
        );

    \I__14470\ : InMux
    port map (
            O => \N__59466\,
            I => \N__59332\
        );

    \I__14469\ : LocalMux
    port map (
            O => \N__59461\,
            I => \N__59317\
        );

    \I__14468\ : LocalMux
    port map (
            O => \N__59458\,
            I => \N__59308\
        );

    \I__14467\ : LocalMux
    port map (
            O => \N__59455\,
            I => \N__59308\
        );

    \I__14466\ : LocalMux
    port map (
            O => \N__59450\,
            I => \N__59308\
        );

    \I__14465\ : LocalMux
    port map (
            O => \N__59447\,
            I => \N__59308\
        );

    \I__14464\ : InMux
    port map (
            O => \N__59446\,
            I => \N__59298\
        );

    \I__14463\ : InMux
    port map (
            O => \N__59445\,
            I => \N__59298\
        );

    \I__14462\ : InMux
    port map (
            O => \N__59444\,
            I => \N__59298\
        );

    \I__14461\ : InMux
    port map (
            O => \N__59443\,
            I => \N__59293\
        );

    \I__14460\ : InMux
    port map (
            O => \N__59442\,
            I => \N__59293\
        );

    \I__14459\ : InMux
    port map (
            O => \N__59441\,
            I => \N__59288\
        );

    \I__14458\ : InMux
    port map (
            O => \N__59440\,
            I => \N__59288\
        );

    \I__14457\ : InMux
    port map (
            O => \N__59439\,
            I => \N__59283\
        );

    \I__14456\ : InMux
    port map (
            O => \N__59438\,
            I => \N__59283\
        );

    \I__14455\ : InMux
    port map (
            O => \N__59437\,
            I => \N__59278\
        );

    \I__14454\ : InMux
    port map (
            O => \N__59436\,
            I => \N__59278\
        );

    \I__14453\ : InMux
    port map (
            O => \N__59435\,
            I => \N__59269\
        );

    \I__14452\ : InMux
    port map (
            O => \N__59434\,
            I => \N__59269\
        );

    \I__14451\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59269\
        );

    \I__14450\ : InMux
    port map (
            O => \N__59432\,
            I => \N__59269\
        );

    \I__14449\ : InMux
    port map (
            O => \N__59431\,
            I => \N__59258\
        );

    \I__14448\ : InMux
    port map (
            O => \N__59430\,
            I => \N__59251\
        );

    \I__14447\ : InMux
    port map (
            O => \N__59429\,
            I => \N__59251\
        );

    \I__14446\ : InMux
    port map (
            O => \N__59428\,
            I => \N__59251\
        );

    \I__14445\ : InMux
    port map (
            O => \N__59427\,
            I => \N__59247\
        );

    \I__14444\ : InMux
    port map (
            O => \N__59426\,
            I => \N__59241\
        );

    \I__14443\ : InMux
    port map (
            O => \N__59425\,
            I => \N__59241\
        );

    \I__14442\ : InMux
    port map (
            O => \N__59424\,
            I => \N__59238\
        );

    \I__14441\ : InMux
    port map (
            O => \N__59423\,
            I => \N__59231\
        );

    \I__14440\ : InMux
    port map (
            O => \N__59422\,
            I => \N__59231\
        );

    \I__14439\ : InMux
    port map (
            O => \N__59421\,
            I => \N__59231\
        );

    \I__14438\ : InMux
    port map (
            O => \N__59420\,
            I => \N__59228\
        );

    \I__14437\ : LocalMux
    port map (
            O => \N__59417\,
            I => \N__59218\
        );

    \I__14436\ : LocalMux
    port map (
            O => \N__59414\,
            I => \N__59218\
        );

    \I__14435\ : LocalMux
    port map (
            O => \N__59411\,
            I => \N__59218\
        );

    \I__14434\ : InMux
    port map (
            O => \N__59410\,
            I => \N__59215\
        );

    \I__14433\ : InMux
    port map (
            O => \N__59409\,
            I => \N__59210\
        );

    \I__14432\ : InMux
    port map (
            O => \N__59408\,
            I => \N__59210\
        );

    \I__14431\ : InMux
    port map (
            O => \N__59407\,
            I => \N__59206\
        );

    \I__14430\ : InMux
    port map (
            O => \N__59406\,
            I => \N__59201\
        );

    \I__14429\ : InMux
    port map (
            O => \N__59405\,
            I => \N__59201\
        );

    \I__14428\ : LocalMux
    port map (
            O => \N__59402\,
            I => \N__59198\
        );

    \I__14427\ : InMux
    port map (
            O => \N__59401\,
            I => \N__59193\
        );

    \I__14426\ : InMux
    port map (
            O => \N__59400\,
            I => \N__59193\
        );

    \I__14425\ : InMux
    port map (
            O => \N__59399\,
            I => \N__59186\
        );

    \I__14424\ : InMux
    port map (
            O => \N__59398\,
            I => \N__59182\
        );

    \I__14423\ : InMux
    port map (
            O => \N__59397\,
            I => \N__59178\
        );

    \I__14422\ : Span4Mux_v
    port map (
            O => \N__59394\,
            I => \N__59165\
        );

    \I__14421\ : LocalMux
    port map (
            O => \N__59391\,
            I => \N__59165\
        );

    \I__14420\ : LocalMux
    port map (
            O => \N__59388\,
            I => \N__59165\
        );

    \I__14419\ : LocalMux
    port map (
            O => \N__59381\,
            I => \N__59165\
        );

    \I__14418\ : Span4Mux_h
    port map (
            O => \N__59378\,
            I => \N__59165\
        );

    \I__14417\ : LocalMux
    port map (
            O => \N__59373\,
            I => \N__59165\
        );

    \I__14416\ : InMux
    port map (
            O => \N__59372\,
            I => \N__59160\
        );

    \I__14415\ : InMux
    port map (
            O => \N__59371\,
            I => \N__59160\
        );

    \I__14414\ : LocalMux
    port map (
            O => \N__59368\,
            I => \N__59157\
        );

    \I__14413\ : InMux
    port map (
            O => \N__59367\,
            I => \N__59148\
        );

    \I__14412\ : InMux
    port map (
            O => \N__59366\,
            I => \N__59148\
        );

    \I__14411\ : InMux
    port map (
            O => \N__59365\,
            I => \N__59148\
        );

    \I__14410\ : InMux
    port map (
            O => \N__59364\,
            I => \N__59148\
        );

    \I__14409\ : InMux
    port map (
            O => \N__59363\,
            I => \N__59143\
        );

    \I__14408\ : InMux
    port map (
            O => \N__59362\,
            I => \N__59143\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__59359\,
            I => \N__59138\
        );

    \I__14406\ : LocalMux
    port map (
            O => \N__59356\,
            I => \N__59138\
        );

    \I__14405\ : InMux
    port map (
            O => \N__59355\,
            I => \N__59127\
        );

    \I__14404\ : InMux
    port map (
            O => \N__59354\,
            I => \N__59127\
        );

    \I__14403\ : InMux
    port map (
            O => \N__59353\,
            I => \N__59127\
        );

    \I__14402\ : InMux
    port map (
            O => \N__59352\,
            I => \N__59127\
        );

    \I__14401\ : InMux
    port map (
            O => \N__59351\,
            I => \N__59127\
        );

    \I__14400\ : InMux
    port map (
            O => \N__59350\,
            I => \N__59124\
        );

    \I__14399\ : LocalMux
    port map (
            O => \N__59347\,
            I => \N__59121\
        );

    \I__14398\ : Span4Mux_v
    port map (
            O => \N__59342\,
            I => \N__59116\
        );

    \I__14397\ : LocalMux
    port map (
            O => \N__59337\,
            I => \N__59116\
        );

    \I__14396\ : InMux
    port map (
            O => \N__59336\,
            I => \N__59106\
        );

    \I__14395\ : InMux
    port map (
            O => \N__59335\,
            I => \N__59106\
        );

    \I__14394\ : LocalMux
    port map (
            O => \N__59332\,
            I => \N__59103\
        );

    \I__14393\ : InMux
    port map (
            O => \N__59331\,
            I => \N__59094\
        );

    \I__14392\ : InMux
    port map (
            O => \N__59330\,
            I => \N__59094\
        );

    \I__14391\ : InMux
    port map (
            O => \N__59329\,
            I => \N__59094\
        );

    \I__14390\ : InMux
    port map (
            O => \N__59328\,
            I => \N__59094\
        );

    \I__14389\ : InMux
    port map (
            O => \N__59327\,
            I => \N__59091\
        );

    \I__14388\ : InMux
    port map (
            O => \N__59326\,
            I => \N__59082\
        );

    \I__14387\ : InMux
    port map (
            O => \N__59325\,
            I => \N__59082\
        );

    \I__14386\ : InMux
    port map (
            O => \N__59324\,
            I => \N__59082\
        );

    \I__14385\ : InMux
    port map (
            O => \N__59323\,
            I => \N__59082\
        );

    \I__14384\ : InMux
    port map (
            O => \N__59322\,
            I => \N__59079\
        );

    \I__14383\ : InMux
    port map (
            O => \N__59321\,
            I => \N__59074\
        );

    \I__14382\ : InMux
    port map (
            O => \N__59320\,
            I => \N__59074\
        );

    \I__14381\ : Span4Mux_v
    port map (
            O => \N__59317\,
            I => \N__59069\
        );

    \I__14380\ : Span4Mux_v
    port map (
            O => \N__59308\,
            I => \N__59069\
        );

    \I__14379\ : InMux
    port map (
            O => \N__59307\,
            I => \N__59066\
        );

    \I__14378\ : InMux
    port map (
            O => \N__59306\,
            I => \N__59063\
        );

    \I__14377\ : InMux
    port map (
            O => \N__59305\,
            I => \N__59060\
        );

    \I__14376\ : LocalMux
    port map (
            O => \N__59298\,
            I => \N__59057\
        );

    \I__14375\ : LocalMux
    port map (
            O => \N__59293\,
            I => \N__59050\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__59288\,
            I => \N__59050\
        );

    \I__14373\ : LocalMux
    port map (
            O => \N__59283\,
            I => \N__59050\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__59278\,
            I => \N__59045\
        );

    \I__14371\ : LocalMux
    port map (
            O => \N__59269\,
            I => \N__59045\
        );

    \I__14370\ : InMux
    port map (
            O => \N__59268\,
            I => \N__59042\
        );

    \I__14369\ : InMux
    port map (
            O => \N__59267\,
            I => \N__59035\
        );

    \I__14368\ : InMux
    port map (
            O => \N__59266\,
            I => \N__59035\
        );

    \I__14367\ : InMux
    port map (
            O => \N__59265\,
            I => \N__59035\
        );

    \I__14366\ : InMux
    port map (
            O => \N__59264\,
            I => \N__59026\
        );

    \I__14365\ : InMux
    port map (
            O => \N__59263\,
            I => \N__59026\
        );

    \I__14364\ : InMux
    port map (
            O => \N__59262\,
            I => \N__59026\
        );

    \I__14363\ : InMux
    port map (
            O => \N__59261\,
            I => \N__59026\
        );

    \I__14362\ : LocalMux
    port map (
            O => \N__59258\,
            I => \N__59021\
        );

    \I__14361\ : LocalMux
    port map (
            O => \N__59251\,
            I => \N__59021\
        );

    \I__14360\ : InMux
    port map (
            O => \N__59250\,
            I => \N__59017\
        );

    \I__14359\ : LocalMux
    port map (
            O => \N__59247\,
            I => \N__59011\
        );

    \I__14358\ : InMux
    port map (
            O => \N__59246\,
            I => \N__59006\
        );

    \I__14357\ : LocalMux
    port map (
            O => \N__59241\,
            I => \N__58999\
        );

    \I__14356\ : LocalMux
    port map (
            O => \N__59238\,
            I => \N__58999\
        );

    \I__14355\ : LocalMux
    port map (
            O => \N__59231\,
            I => \N__58999\
        );

    \I__14354\ : LocalMux
    port map (
            O => \N__59228\,
            I => \N__58996\
        );

    \I__14353\ : InMux
    port map (
            O => \N__59227\,
            I => \N__58993\
        );

    \I__14352\ : InMux
    port map (
            O => \N__59226\,
            I => \N__58988\
        );

    \I__14351\ : InMux
    port map (
            O => \N__59225\,
            I => \N__58988\
        );

    \I__14350\ : Span4Mux_v
    port map (
            O => \N__59218\,
            I => \N__58981\
        );

    \I__14349\ : LocalMux
    port map (
            O => \N__59215\,
            I => \N__58981\
        );

    \I__14348\ : LocalMux
    port map (
            O => \N__59210\,
            I => \N__58981\
        );

    \I__14347\ : InMux
    port map (
            O => \N__59209\,
            I => \N__58978\
        );

    \I__14346\ : LocalMux
    port map (
            O => \N__59206\,
            I => \N__58973\
        );

    \I__14345\ : LocalMux
    port map (
            O => \N__59201\,
            I => \N__58973\
        );

    \I__14344\ : Span4Mux_v
    port map (
            O => \N__59198\,
            I => \N__58968\
        );

    \I__14343\ : LocalMux
    port map (
            O => \N__59193\,
            I => \N__58968\
        );

    \I__14342\ : InMux
    port map (
            O => \N__59192\,
            I => \N__58963\
        );

    \I__14341\ : InMux
    port map (
            O => \N__59191\,
            I => \N__58963\
        );

    \I__14340\ : InMux
    port map (
            O => \N__59190\,
            I => \N__58960\
        );

    \I__14339\ : InMux
    port map (
            O => \N__59189\,
            I => \N__58957\
        );

    \I__14338\ : LocalMux
    port map (
            O => \N__59186\,
            I => \N__58954\
        );

    \I__14337\ : InMux
    port map (
            O => \N__59185\,
            I => \N__58951\
        );

    \I__14336\ : LocalMux
    port map (
            O => \N__59182\,
            I => \N__58945\
        );

    \I__14335\ : InMux
    port map (
            O => \N__59181\,
            I => \N__58942\
        );

    \I__14334\ : LocalMux
    port map (
            O => \N__59178\,
            I => \N__58939\
        );

    \I__14333\ : Span4Mux_v
    port map (
            O => \N__59165\,
            I => \N__58934\
        );

    \I__14332\ : LocalMux
    port map (
            O => \N__59160\,
            I => \N__58934\
        );

    \I__14331\ : Span4Mux_v
    port map (
            O => \N__59157\,
            I => \N__58923\
        );

    \I__14330\ : LocalMux
    port map (
            O => \N__59148\,
            I => \N__58923\
        );

    \I__14329\ : LocalMux
    port map (
            O => \N__59143\,
            I => \N__58923\
        );

    \I__14328\ : Span4Mux_v
    port map (
            O => \N__59138\,
            I => \N__58923\
        );

    \I__14327\ : LocalMux
    port map (
            O => \N__59127\,
            I => \N__58923\
        );

    \I__14326\ : LocalMux
    port map (
            O => \N__59124\,
            I => \N__58916\
        );

    \I__14325\ : Span4Mux_h
    port map (
            O => \N__59121\,
            I => \N__58916\
        );

    \I__14324\ : Span4Mux_h
    port map (
            O => \N__59116\,
            I => \N__58916\
        );

    \I__14323\ : InMux
    port map (
            O => \N__59115\,
            I => \N__58908\
        );

    \I__14322\ : InMux
    port map (
            O => \N__59114\,
            I => \N__58908\
        );

    \I__14321\ : InMux
    port map (
            O => \N__59113\,
            I => \N__58908\
        );

    \I__14320\ : InMux
    port map (
            O => \N__59112\,
            I => \N__58905\
        );

    \I__14319\ : InMux
    port map (
            O => \N__59111\,
            I => \N__58902\
        );

    \I__14318\ : LocalMux
    port map (
            O => \N__59106\,
            I => \N__58899\
        );

    \I__14317\ : Span4Mux_v
    port map (
            O => \N__59103\,
            I => \N__58896\
        );

    \I__14316\ : LocalMux
    port map (
            O => \N__59094\,
            I => \N__58889\
        );

    \I__14315\ : LocalMux
    port map (
            O => \N__59091\,
            I => \N__58889\
        );

    \I__14314\ : LocalMux
    port map (
            O => \N__59082\,
            I => \N__58889\
        );

    \I__14313\ : LocalMux
    port map (
            O => \N__59079\,
            I => \N__58870\
        );

    \I__14312\ : LocalMux
    port map (
            O => \N__59074\,
            I => \N__58870\
        );

    \I__14311\ : Span4Mux_h
    port map (
            O => \N__59069\,
            I => \N__58870\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__59066\,
            I => \N__58870\
        );

    \I__14309\ : LocalMux
    port map (
            O => \N__59063\,
            I => \N__58870\
        );

    \I__14308\ : LocalMux
    port map (
            O => \N__59060\,
            I => \N__58870\
        );

    \I__14307\ : Span4Mux_h
    port map (
            O => \N__59057\,
            I => \N__58870\
        );

    \I__14306\ : Span4Mux_v
    port map (
            O => \N__59050\,
            I => \N__58870\
        );

    \I__14305\ : Span4Mux_v
    port map (
            O => \N__59045\,
            I => \N__58870\
        );

    \I__14304\ : LocalMux
    port map (
            O => \N__59042\,
            I => \N__58861\
        );

    \I__14303\ : LocalMux
    port map (
            O => \N__59035\,
            I => \N__58861\
        );

    \I__14302\ : LocalMux
    port map (
            O => \N__59026\,
            I => \N__58861\
        );

    \I__14301\ : Span4Mux_v
    port map (
            O => \N__59021\,
            I => \N__58861\
        );

    \I__14300\ : InMux
    port map (
            O => \N__59020\,
            I => \N__58858\
        );

    \I__14299\ : LocalMux
    port map (
            O => \N__59017\,
            I => \N__58852\
        );

    \I__14298\ : InMux
    port map (
            O => \N__59016\,
            I => \N__58845\
        );

    \I__14297\ : InMux
    port map (
            O => \N__59015\,
            I => \N__58845\
        );

    \I__14296\ : InMux
    port map (
            O => \N__59014\,
            I => \N__58845\
        );

    \I__14295\ : Span4Mux_h
    port map (
            O => \N__59011\,
            I => \N__58837\
        );

    \I__14294\ : InMux
    port map (
            O => \N__59010\,
            I => \N__58831\
        );

    \I__14293\ : InMux
    port map (
            O => \N__59009\,
            I => \N__58831\
        );

    \I__14292\ : LocalMux
    port map (
            O => \N__59006\,
            I => \N__58828\
        );

    \I__14291\ : Span4Mux_v
    port map (
            O => \N__58999\,
            I => \N__58823\
        );

    \I__14290\ : Span4Mux_v
    port map (
            O => \N__58996\,
            I => \N__58823\
        );

    \I__14289\ : LocalMux
    port map (
            O => \N__58993\,
            I => \N__58814\
        );

    \I__14288\ : LocalMux
    port map (
            O => \N__58988\,
            I => \N__58814\
        );

    \I__14287\ : Span4Mux_h
    port map (
            O => \N__58981\,
            I => \N__58814\
        );

    \I__14286\ : LocalMux
    port map (
            O => \N__58978\,
            I => \N__58814\
        );

    \I__14285\ : Span4Mux_v
    port map (
            O => \N__58973\,
            I => \N__58807\
        );

    \I__14284\ : Span4Mux_v
    port map (
            O => \N__58968\,
            I => \N__58807\
        );

    \I__14283\ : LocalMux
    port map (
            O => \N__58963\,
            I => \N__58807\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__58960\,
            I => \N__58798\
        );

    \I__14281\ : LocalMux
    port map (
            O => \N__58957\,
            I => \N__58798\
        );

    \I__14280\ : Span4Mux_h
    port map (
            O => \N__58954\,
            I => \N__58798\
        );

    \I__14279\ : LocalMux
    port map (
            O => \N__58951\,
            I => \N__58798\
        );

    \I__14278\ : InMux
    port map (
            O => \N__58950\,
            I => \N__58791\
        );

    \I__14277\ : InMux
    port map (
            O => \N__58949\,
            I => \N__58791\
        );

    \I__14276\ : InMux
    port map (
            O => \N__58948\,
            I => \N__58791\
        );

    \I__14275\ : Span4Mux_h
    port map (
            O => \N__58945\,
            I => \N__58784\
        );

    \I__14274\ : LocalMux
    port map (
            O => \N__58942\,
            I => \N__58784\
        );

    \I__14273\ : Span4Mux_v
    port map (
            O => \N__58939\,
            I => \N__58784\
        );

    \I__14272\ : Span4Mux_h
    port map (
            O => \N__58934\,
            I => \N__58777\
        );

    \I__14271\ : Span4Mux_v
    port map (
            O => \N__58923\,
            I => \N__58777\
        );

    \I__14270\ : Span4Mux_h
    port map (
            O => \N__58916\,
            I => \N__58777\
        );

    \I__14269\ : InMux
    port map (
            O => \N__58915\,
            I => \N__58774\
        );

    \I__14268\ : LocalMux
    port map (
            O => \N__58908\,
            I => \N__58771\
        );

    \I__14267\ : LocalMux
    port map (
            O => \N__58905\,
            I => \N__58766\
        );

    \I__14266\ : LocalMux
    port map (
            O => \N__58902\,
            I => \N__58766\
        );

    \I__14265\ : Span4Mux_h
    port map (
            O => \N__58899\,
            I => \N__58753\
        );

    \I__14264\ : Span4Mux_h
    port map (
            O => \N__58896\,
            I => \N__58753\
        );

    \I__14263\ : Span4Mux_v
    port map (
            O => \N__58889\,
            I => \N__58753\
        );

    \I__14262\ : Span4Mux_v
    port map (
            O => \N__58870\,
            I => \N__58753\
        );

    \I__14261\ : Span4Mux_v
    port map (
            O => \N__58861\,
            I => \N__58753\
        );

    \I__14260\ : LocalMux
    port map (
            O => \N__58858\,
            I => \N__58753\
        );

    \I__14259\ : InMux
    port map (
            O => \N__58857\,
            I => \N__58746\
        );

    \I__14258\ : InMux
    port map (
            O => \N__58856\,
            I => \N__58746\
        );

    \I__14257\ : InMux
    port map (
            O => \N__58855\,
            I => \N__58746\
        );

    \I__14256\ : Span4Mux_h
    port map (
            O => \N__58852\,
            I => \N__58743\
        );

    \I__14255\ : LocalMux
    port map (
            O => \N__58845\,
            I => \N__58740\
        );

    \I__14254\ : InMux
    port map (
            O => \N__58844\,
            I => \N__58733\
        );

    \I__14253\ : InMux
    port map (
            O => \N__58843\,
            I => \N__58733\
        );

    \I__14252\ : InMux
    port map (
            O => \N__58842\,
            I => \N__58733\
        );

    \I__14251\ : InMux
    port map (
            O => \N__58841\,
            I => \N__58730\
        );

    \I__14250\ : InMux
    port map (
            O => \N__58840\,
            I => \N__58727\
        );

    \I__14249\ : Span4Mux_v
    port map (
            O => \N__58837\,
            I => \N__58724\
        );

    \I__14248\ : InMux
    port map (
            O => \N__58836\,
            I => \N__58721\
        );

    \I__14247\ : LocalMux
    port map (
            O => \N__58831\,
            I => \N__58716\
        );

    \I__14246\ : Span12Mux_h
    port map (
            O => \N__58828\,
            I => \N__58716\
        );

    \I__14245\ : Span4Mux_h
    port map (
            O => \N__58823\,
            I => \N__58709\
        );

    \I__14244\ : Span4Mux_v
    port map (
            O => \N__58814\,
            I => \N__58709\
        );

    \I__14243\ : Span4Mux_h
    port map (
            O => \N__58807\,
            I => \N__58709\
        );

    \I__14242\ : Span4Mux_v
    port map (
            O => \N__58798\,
            I => \N__58700\
        );

    \I__14241\ : LocalMux
    port map (
            O => \N__58791\,
            I => \N__58700\
        );

    \I__14240\ : Span4Mux_h
    port map (
            O => \N__58784\,
            I => \N__58700\
        );

    \I__14239\ : Span4Mux_h
    port map (
            O => \N__58777\,
            I => \N__58700\
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__58774\,
            I => \N__58689\
        );

    \I__14237\ : Span12Mux_v
    port map (
            O => \N__58771\,
            I => \N__58689\
        );

    \I__14236\ : Span12Mux_h
    port map (
            O => \N__58766\,
            I => \N__58689\
        );

    \I__14235\ : Sp12to4
    port map (
            O => \N__58753\,
            I => \N__58689\
        );

    \I__14234\ : LocalMux
    port map (
            O => \N__58746\,
            I => \N__58689\
        );

    \I__14233\ : Odrv4
    port map (
            O => \N__58743\,
            I => comm_cmd_0
        );

    \I__14232\ : Odrv4
    port map (
            O => \N__58740\,
            I => comm_cmd_0
        );

    \I__14231\ : LocalMux
    port map (
            O => \N__58733\,
            I => comm_cmd_0
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__58730\,
            I => comm_cmd_0
        );

    \I__14229\ : LocalMux
    port map (
            O => \N__58727\,
            I => comm_cmd_0
        );

    \I__14228\ : Odrv4
    port map (
            O => \N__58724\,
            I => comm_cmd_0
        );

    \I__14227\ : LocalMux
    port map (
            O => \N__58721\,
            I => comm_cmd_0
        );

    \I__14226\ : Odrv12
    port map (
            O => \N__58716\,
            I => comm_cmd_0
        );

    \I__14225\ : Odrv4
    port map (
            O => \N__58709\,
            I => comm_cmd_0
        );

    \I__14224\ : Odrv4
    port map (
            O => \N__58700\,
            I => comm_cmd_0
        );

    \I__14223\ : Odrv12
    port map (
            O => \N__58689\,
            I => comm_cmd_0
        );

    \I__14222\ : InMux
    port map (
            O => \N__58666\,
            I => \N__58663\
        );

    \I__14221\ : LocalMux
    port map (
            O => \N__58663\,
            I => \N__58660\
        );

    \I__14220\ : Span4Mux_h
    port map (
            O => \N__58660\,
            I => \N__58657\
        );

    \I__14219\ : Odrv4
    port map (
            O => \N__58657\,
            I => n22649
        );

    \I__14218\ : InMux
    port map (
            O => \N__58654\,
            I => \N__58643\
        );

    \I__14217\ : InMux
    port map (
            O => \N__58653\,
            I => \N__58643\
        );

    \I__14216\ : InMux
    port map (
            O => \N__58652\,
            I => \N__58638\
        );

    \I__14215\ : InMux
    port map (
            O => \N__58651\,
            I => \N__58635\
        );

    \I__14214\ : InMux
    port map (
            O => \N__58650\,
            I => \N__58630\
        );

    \I__14213\ : InMux
    port map (
            O => \N__58649\,
            I => \N__58630\
        );

    \I__14212\ : InMux
    port map (
            O => \N__58648\,
            I => \N__58627\
        );

    \I__14211\ : LocalMux
    port map (
            O => \N__58643\,
            I => \N__58621\
        );

    \I__14210\ : InMux
    port map (
            O => \N__58642\,
            I => \N__58616\
        );

    \I__14209\ : InMux
    port map (
            O => \N__58641\,
            I => \N__58616\
        );

    \I__14208\ : LocalMux
    port map (
            O => \N__58638\,
            I => \N__58611\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__58635\,
            I => \N__58602\
        );

    \I__14206\ : LocalMux
    port map (
            O => \N__58630\,
            I => \N__58602\
        );

    \I__14205\ : LocalMux
    port map (
            O => \N__58627\,
            I => \N__58599\
        );

    \I__14204\ : InMux
    port map (
            O => \N__58626\,
            I => \N__58594\
        );

    \I__14203\ : InMux
    port map (
            O => \N__58625\,
            I => \N__58594\
        );

    \I__14202\ : InMux
    port map (
            O => \N__58624\,
            I => \N__58591\
        );

    \I__14201\ : Span4Mux_v
    port map (
            O => \N__58621\,
            I => \N__58586\
        );

    \I__14200\ : LocalMux
    port map (
            O => \N__58616\,
            I => \N__58586\
        );

    \I__14199\ : InMux
    port map (
            O => \N__58615\,
            I => \N__58581\
        );

    \I__14198\ : InMux
    port map (
            O => \N__58614\,
            I => \N__58578\
        );

    \I__14197\ : Span4Mux_h
    port map (
            O => \N__58611\,
            I => \N__58575\
        );

    \I__14196\ : InMux
    port map (
            O => \N__58610\,
            I => \N__58572\
        );

    \I__14195\ : InMux
    port map (
            O => \N__58609\,
            I => \N__58567\
        );

    \I__14194\ : InMux
    port map (
            O => \N__58608\,
            I => \N__58567\
        );

    \I__14193\ : InMux
    port map (
            O => \N__58607\,
            I => \N__58564\
        );

    \I__14192\ : Span4Mux_v
    port map (
            O => \N__58602\,
            I => \N__58557\
        );

    \I__14191\ : Span4Mux_v
    port map (
            O => \N__58599\,
            I => \N__58557\
        );

    \I__14190\ : LocalMux
    port map (
            O => \N__58594\,
            I => \N__58557\
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__58591\,
            I => \N__58552\
        );

    \I__14188\ : Span4Mux_h
    port map (
            O => \N__58586\,
            I => \N__58552\
        );

    \I__14187\ : InMux
    port map (
            O => \N__58585\,
            I => \N__58547\
        );

    \I__14186\ : InMux
    port map (
            O => \N__58584\,
            I => \N__58547\
        );

    \I__14185\ : LocalMux
    port map (
            O => \N__58581\,
            I => comm_cmd_5
        );

    \I__14184\ : LocalMux
    port map (
            O => \N__58578\,
            I => comm_cmd_5
        );

    \I__14183\ : Odrv4
    port map (
            O => \N__58575\,
            I => comm_cmd_5
        );

    \I__14182\ : LocalMux
    port map (
            O => \N__58572\,
            I => comm_cmd_5
        );

    \I__14181\ : LocalMux
    port map (
            O => \N__58567\,
            I => comm_cmd_5
        );

    \I__14180\ : LocalMux
    port map (
            O => \N__58564\,
            I => comm_cmd_5
        );

    \I__14179\ : Odrv4
    port map (
            O => \N__58557\,
            I => comm_cmd_5
        );

    \I__14178\ : Odrv4
    port map (
            O => \N__58552\,
            I => comm_cmd_5
        );

    \I__14177\ : LocalMux
    port map (
            O => \N__58547\,
            I => comm_cmd_5
        );

    \I__14176\ : InMux
    port map (
            O => \N__58528\,
            I => \N__58523\
        );

    \I__14175\ : InMux
    port map (
            O => \N__58527\,
            I => \N__58516\
        );

    \I__14174\ : InMux
    port map (
            O => \N__58526\,
            I => \N__58516\
        );

    \I__14173\ : LocalMux
    port map (
            O => \N__58523\,
            I => \N__58512\
        );

    \I__14172\ : InMux
    port map (
            O => \N__58522\,
            I => \N__58508\
        );

    \I__14171\ : CascadeMux
    port map (
            O => \N__58521\,
            I => \N__58505\
        );

    \I__14170\ : LocalMux
    port map (
            O => \N__58516\,
            I => \N__58502\
        );

    \I__14169\ : InMux
    port map (
            O => \N__58515\,
            I => \N__58499\
        );

    \I__14168\ : Span4Mux_v
    port map (
            O => \N__58512\,
            I => \N__58496\
        );

    \I__14167\ : CascadeMux
    port map (
            O => \N__58511\,
            I => \N__58493\
        );

    \I__14166\ : LocalMux
    port map (
            O => \N__58508\,
            I => \N__58488\
        );

    \I__14165\ : InMux
    port map (
            O => \N__58505\,
            I => \N__58484\
        );

    \I__14164\ : Span4Mux_v
    port map (
            O => \N__58502\,
            I => \N__58475\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__58499\,
            I => \N__58475\
        );

    \I__14162\ : Span4Mux_v
    port map (
            O => \N__58496\,
            I => \N__58475\
        );

    \I__14161\ : InMux
    port map (
            O => \N__58493\,
            I => \N__58470\
        );

    \I__14160\ : InMux
    port map (
            O => \N__58492\,
            I => \N__58470\
        );

    \I__14159\ : CascadeMux
    port map (
            O => \N__58491\,
            I => \N__58466\
        );

    \I__14158\ : Span4Mux_h
    port map (
            O => \N__58488\,
            I => \N__58463\
        );

    \I__14157\ : InMux
    port map (
            O => \N__58487\,
            I => \N__58460\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__58484\,
            I => \N__58457\
        );

    \I__14155\ : InMux
    port map (
            O => \N__58483\,
            I => \N__58452\
        );

    \I__14154\ : InMux
    port map (
            O => \N__58482\,
            I => \N__58452\
        );

    \I__14153\ : Sp12to4
    port map (
            O => \N__58475\,
            I => \N__58447\
        );

    \I__14152\ : LocalMux
    port map (
            O => \N__58470\,
            I => \N__58447\
        );

    \I__14151\ : InMux
    port map (
            O => \N__58469\,
            I => \N__58442\
        );

    \I__14150\ : InMux
    port map (
            O => \N__58466\,
            I => \N__58442\
        );

    \I__14149\ : Odrv4
    port map (
            O => \N__58463\,
            I => comm_cmd_4
        );

    \I__14148\ : LocalMux
    port map (
            O => \N__58460\,
            I => comm_cmd_4
        );

    \I__14147\ : Odrv4
    port map (
            O => \N__58457\,
            I => comm_cmd_4
        );

    \I__14146\ : LocalMux
    port map (
            O => \N__58452\,
            I => comm_cmd_4
        );

    \I__14145\ : Odrv12
    port map (
            O => \N__58447\,
            I => comm_cmd_4
        );

    \I__14144\ : LocalMux
    port map (
            O => \N__58442\,
            I => comm_cmd_4
        );

    \I__14143\ : InMux
    port map (
            O => \N__58429\,
            I => \N__58426\
        );

    \I__14142\ : LocalMux
    port map (
            O => \N__58426\,
            I => n22365
        );

    \I__14141\ : CascadeMux
    port map (
            O => \N__58423\,
            I => \n22364_cascade_\
        );

    \I__14140\ : InMux
    port map (
            O => \N__58420\,
            I => \N__58417\
        );

    \I__14139\ : LocalMux
    port map (
            O => \N__58417\,
            I => n48
        );

    \I__14138\ : CascadeMux
    port map (
            O => \N__58414\,
            I => \n22370_cascade_\
        );

    \I__14137\ : InMux
    port map (
            O => \N__58411\,
            I => \N__58408\
        );

    \I__14136\ : LocalMux
    port map (
            O => \N__58408\,
            I => \N__58404\
        );

    \I__14135\ : InMux
    port map (
            O => \N__58407\,
            I => \N__58400\
        );

    \I__14134\ : Span4Mux_h
    port map (
            O => \N__58404\,
            I => \N__58396\
        );

    \I__14133\ : InMux
    port map (
            O => \N__58403\,
            I => \N__58393\
        );

    \I__14132\ : LocalMux
    port map (
            O => \N__58400\,
            I => \N__58390\
        );

    \I__14131\ : InMux
    port map (
            O => \N__58399\,
            I => \N__58387\
        );

    \I__14130\ : Odrv4
    port map (
            O => \N__58396\,
            I => n7148
        );

    \I__14129\ : LocalMux
    port map (
            O => \N__58393\,
            I => n7148
        );

    \I__14128\ : Odrv4
    port map (
            O => \N__58390\,
            I => n7148
        );

    \I__14127\ : LocalMux
    port map (
            O => \N__58387\,
            I => n7148
        );

    \I__14126\ : InMux
    port map (
            O => \N__58378\,
            I => \N__58375\
        );

    \I__14125\ : LocalMux
    port map (
            O => \N__58375\,
            I => \N__58372\
        );

    \I__14124\ : Odrv4
    port map (
            O => \N__58372\,
            I => n22368
        );

    \I__14123\ : InMux
    port map (
            O => \N__58369\,
            I => \N__58366\
        );

    \I__14122\ : LocalMux
    port map (
            O => \N__58366\,
            I => \N__58362\
        );

    \I__14121\ : InMux
    port map (
            O => \N__58365\,
            I => \N__58359\
        );

    \I__14120\ : Span4Mux_h
    port map (
            O => \N__58362\,
            I => \N__58356\
        );

    \I__14119\ : LocalMux
    port map (
            O => \N__58359\,
            I => \N__58353\
        );

    \I__14118\ : Odrv4
    port map (
            O => \N__58356\,
            I => n9_adj_1507
        );

    \I__14117\ : Odrv12
    port map (
            O => \N__58353\,
            I => n9_adj_1507
        );

    \I__14116\ : InMux
    port map (
            O => \N__58348\,
            I => \N__58345\
        );

    \I__14115\ : LocalMux
    port map (
            O => \N__58345\,
            I => \N__58342\
        );

    \I__14114\ : Span4Mux_v
    port map (
            O => \N__58342\,
            I => \N__58339\
        );

    \I__14113\ : Span4Mux_h
    port map (
            O => \N__58339\,
            I => \N__58336\
        );

    \I__14112\ : Span4Mux_h
    port map (
            O => \N__58336\,
            I => \N__58333\
        );

    \I__14111\ : Odrv4
    port map (
            O => \N__58333\,
            I => n23387
        );

    \I__14110\ : CascadeMux
    port map (
            O => \N__58330\,
            I => \N__58327\
        );

    \I__14109\ : InMux
    port map (
            O => \N__58327\,
            I => \N__58324\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__58324\,
            I => \N__58321\
        );

    \I__14107\ : Odrv4
    port map (
            O => \N__58321\,
            I => n23351
        );

    \I__14106\ : InMux
    port map (
            O => \N__58318\,
            I => \N__58315\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__58315\,
            I => n23495
        );

    \I__14104\ : InMux
    port map (
            O => \N__58312\,
            I => \N__58309\
        );

    \I__14103\ : LocalMux
    port map (
            O => \N__58309\,
            I => \N__58306\
        );

    \I__14102\ : Span4Mux_v
    port map (
            O => \N__58306\,
            I => \N__58303\
        );

    \I__14101\ : Odrv4
    port map (
            O => \N__58303\,
            I => buf_data_iac_19
        );

    \I__14100\ : InMux
    port map (
            O => \N__58300\,
            I => \N__58297\
        );

    \I__14099\ : LocalMux
    port map (
            O => \N__58297\,
            I => \N__58294\
        );

    \I__14098\ : Odrv12
    port map (
            O => \N__58294\,
            I => n22642
        );

    \I__14097\ : CascadeMux
    port map (
            O => \N__58291\,
            I => \N__58288\
        );

    \I__14096\ : InMux
    port map (
            O => \N__58288\,
            I => \N__58285\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__58285\,
            I => \N__58282\
        );

    \I__14094\ : Span4Mux_h
    port map (
            O => \N__58282\,
            I => \N__58279\
        );

    \I__14093\ : Odrv4
    port map (
            O => \N__58279\,
            I => n23_adj_1791
        );

    \I__14092\ : InMux
    port map (
            O => \N__58276\,
            I => \N__58273\
        );

    \I__14091\ : LocalMux
    port map (
            O => \N__58273\,
            I => \N__58270\
        );

    \I__14090\ : Span4Mux_v
    port map (
            O => \N__58270\,
            I => \N__58267\
        );

    \I__14089\ : Sp12to4
    port map (
            O => \N__58267\,
            I => \N__58264\
        );

    \I__14088\ : Span12Mux_h
    port map (
            O => \N__58264\,
            I => \N__58261\
        );

    \I__14087\ : Odrv12
    port map (
            O => \N__58261\,
            I => n23501
        );

    \I__14086\ : CascadeMux
    port map (
            O => \N__58258\,
            I => \n23459_cascade_\
        );

    \I__14085\ : InMux
    port map (
            O => \N__58255\,
            I => \N__58252\
        );

    \I__14084\ : LocalMux
    port map (
            O => \N__58252\,
            I => \N__58249\
        );

    \I__14083\ : Span4Mux_v
    port map (
            O => \N__58249\,
            I => \N__58246\
        );

    \I__14082\ : Sp12to4
    port map (
            O => \N__58246\,
            I => \N__58243\
        );

    \I__14081\ : Span12Mux_h
    port map (
            O => \N__58243\,
            I => \N__58240\
        );

    \I__14080\ : Odrv12
    port map (
            O => \N__58240\,
            I => n112_adj_1795
        );

    \I__14079\ : InMux
    port map (
            O => \N__58237\,
            I => \N__58234\
        );

    \I__14078\ : LocalMux
    port map (
            O => \N__58234\,
            I => n22492
        );

    \I__14077\ : CascadeMux
    port map (
            O => \N__58231\,
            I => \n6_adj_1657_cascade_\
        );

    \I__14076\ : CascadeMux
    port map (
            O => \N__58228\,
            I => \n26_adj_1597_cascade_\
        );

    \I__14075\ : CEMux
    port map (
            O => \N__58225\,
            I => \N__58222\
        );

    \I__14074\ : LocalMux
    port map (
            O => \N__58222\,
            I => \N__58219\
        );

    \I__14073\ : Odrv4
    port map (
            O => \N__58219\,
            I => n18_adj_1595
        );

    \I__14072\ : InMux
    port map (
            O => \N__58216\,
            I => \N__58213\
        );

    \I__14071\ : LocalMux
    port map (
            O => \N__58213\,
            I => n21908
        );

    \I__14070\ : InMux
    port map (
            O => \N__58210\,
            I => \N__58201\
        );

    \I__14069\ : InMux
    port map (
            O => \N__58209\,
            I => \N__58194\
        );

    \I__14068\ : InMux
    port map (
            O => \N__58208\,
            I => \N__58194\
        );

    \I__14067\ : InMux
    port map (
            O => \N__58207\,
            I => \N__58194\
        );

    \I__14066\ : CascadeMux
    port map (
            O => \N__58206\,
            I => \N__58189\
        );

    \I__14065\ : CascadeMux
    port map (
            O => \N__58205\,
            I => \N__58182\
        );

    \I__14064\ : InMux
    port map (
            O => \N__58204\,
            I => \N__58178\
        );

    \I__14063\ : LocalMux
    port map (
            O => \N__58201\,
            I => \N__58173\
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__58194\,
            I => \N__58173\
        );

    \I__14061\ : InMux
    port map (
            O => \N__58193\,
            I => \N__58170\
        );

    \I__14060\ : InMux
    port map (
            O => \N__58192\,
            I => \N__58161\
        );

    \I__14059\ : InMux
    port map (
            O => \N__58189\,
            I => \N__58161\
        );

    \I__14058\ : InMux
    port map (
            O => \N__58188\,
            I => \N__58161\
        );

    \I__14057\ : InMux
    port map (
            O => \N__58187\,
            I => \N__58161\
        );

    \I__14056\ : InMux
    port map (
            O => \N__58186\,
            I => \N__58154\
        );

    \I__14055\ : InMux
    port map (
            O => \N__58185\,
            I => \N__58154\
        );

    \I__14054\ : InMux
    port map (
            O => \N__58182\,
            I => \N__58154\
        );

    \I__14053\ : CascadeMux
    port map (
            O => \N__58181\,
            I => \N__58148\
        );

    \I__14052\ : LocalMux
    port map (
            O => \N__58178\,
            I => \N__58144\
        );

    \I__14051\ : Span4Mux_v
    port map (
            O => \N__58173\,
            I => \N__58141\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__58170\,
            I => \N__58138\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__58161\,
            I => \N__58133\
        );

    \I__14048\ : LocalMux
    port map (
            O => \N__58154\,
            I => \N__58133\
        );

    \I__14047\ : InMux
    port map (
            O => \N__58153\,
            I => \N__58129\
        );

    \I__14046\ : InMux
    port map (
            O => \N__58152\,
            I => \N__58126\
        );

    \I__14045\ : InMux
    port map (
            O => \N__58151\,
            I => \N__58119\
        );

    \I__14044\ : InMux
    port map (
            O => \N__58148\,
            I => \N__58119\
        );

    \I__14043\ : InMux
    port map (
            O => \N__58147\,
            I => \N__58119\
        );

    \I__14042\ : Span4Mux_v
    port map (
            O => \N__58144\,
            I => \N__58114\
        );

    \I__14041\ : Span4Mux_h
    port map (
            O => \N__58141\,
            I => \N__58107\
        );

    \I__14040\ : Span4Mux_h
    port map (
            O => \N__58138\,
            I => \N__58107\
        );

    \I__14039\ : Span4Mux_v
    port map (
            O => \N__58133\,
            I => \N__58107\
        );

    \I__14038\ : CascadeMux
    port map (
            O => \N__58132\,
            I => \N__58104\
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__58129\,
            I => \N__58097\
        );

    \I__14036\ : LocalMux
    port map (
            O => \N__58126\,
            I => \N__58097\
        );

    \I__14035\ : LocalMux
    port map (
            O => \N__58119\,
            I => \N__58097\
        );

    \I__14034\ : InMux
    port map (
            O => \N__58118\,
            I => \N__58092\
        );

    \I__14033\ : InMux
    port map (
            O => \N__58117\,
            I => \N__58092\
        );

    \I__14032\ : Span4Mux_v
    port map (
            O => \N__58114\,
            I => \N__58089\
        );

    \I__14031\ : Span4Mux_h
    port map (
            O => \N__58107\,
            I => \N__58086\
        );

    \I__14030\ : InMux
    port map (
            O => \N__58104\,
            I => \N__58083\
        );

    \I__14029\ : Span4Mux_v
    port map (
            O => \N__58097\,
            I => \N__58080\
        );

    \I__14028\ : LocalMux
    port map (
            O => \N__58092\,
            I => \N__58077\
        );

    \I__14027\ : Span4Mux_v
    port map (
            O => \N__58089\,
            I => \N__58074\
        );

    \I__14026\ : Sp12to4
    port map (
            O => \N__58086\,
            I => \N__58071\
        );

    \I__14025\ : LocalMux
    port map (
            O => \N__58083\,
            I => \N__58068\
        );

    \I__14024\ : Sp12to4
    port map (
            O => \N__58080\,
            I => \N__58063\
        );

    \I__14023\ : Span12Mux_v
    port map (
            O => \N__58077\,
            I => \N__58063\
        );

    \I__14022\ : Sp12to4
    port map (
            O => \N__58074\,
            I => \N__58060\
        );

    \I__14021\ : Span12Mux_s2_h
    port map (
            O => \N__58071\,
            I => \N__58055\
        );

    \I__14020\ : Span12Mux_h
    port map (
            O => \N__58068\,
            I => \N__58055\
        );

    \I__14019\ : Span12Mux_v
    port map (
            O => \N__58063\,
            I => \N__58052\
        );

    \I__14018\ : Span12Mux_h
    port map (
            O => \N__58060\,
            I => \N__58047\
        );

    \I__14017\ : Span12Mux_v
    port map (
            O => \N__58055\,
            I => \N__58047\
        );

    \I__14016\ : Odrv12
    port map (
            O => \N__58052\,
            I => \ICE_SPI_CE0\
        );

    \I__14015\ : Odrv12
    port map (
            O => \N__58047\,
            I => \ICE_SPI_CE0\
        );

    \I__14014\ : InMux
    port map (
            O => \N__58042\,
            I => \N__58023\
        );

    \I__14013\ : InMux
    port map (
            O => \N__58041\,
            I => \N__58023\
        );

    \I__14012\ : InMux
    port map (
            O => \N__58040\,
            I => \N__58023\
        );

    \I__14011\ : CascadeMux
    port map (
            O => \N__58039\,
            I => \N__58019\
        );

    \I__14010\ : InMux
    port map (
            O => \N__58038\,
            I => \N__58011\
        );

    \I__14009\ : InMux
    port map (
            O => \N__58037\,
            I => \N__58011\
        );

    \I__14008\ : InMux
    port map (
            O => \N__58036\,
            I => \N__58011\
        );

    \I__14007\ : InMux
    port map (
            O => \N__58035\,
            I => \N__58002\
        );

    \I__14006\ : InMux
    port map (
            O => \N__58034\,
            I => \N__58002\
        );

    \I__14005\ : InMux
    port map (
            O => \N__58033\,
            I => \N__58002\
        );

    \I__14004\ : InMux
    port map (
            O => \N__58032\,
            I => \N__58002\
        );

    \I__14003\ : InMux
    port map (
            O => \N__58031\,
            I => \N__57999\
        );

    \I__14002\ : InMux
    port map (
            O => \N__58030\,
            I => \N__57996\
        );

    \I__14001\ : LocalMux
    port map (
            O => \N__58023\,
            I => \N__57993\
        );

    \I__14000\ : InMux
    port map (
            O => \N__58022\,
            I => \N__57990\
        );

    \I__13999\ : InMux
    port map (
            O => \N__58019\,
            I => \N__57985\
        );

    \I__13998\ : InMux
    port map (
            O => \N__58018\,
            I => \N__57985\
        );

    \I__13997\ : LocalMux
    port map (
            O => \N__58011\,
            I => comm_data_vld
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__58002\,
            I => comm_data_vld
        );

    \I__13995\ : LocalMux
    port map (
            O => \N__57999\,
            I => comm_data_vld
        );

    \I__13994\ : LocalMux
    port map (
            O => \N__57996\,
            I => comm_data_vld
        );

    \I__13993\ : Odrv4
    port map (
            O => \N__57993\,
            I => comm_data_vld
        );

    \I__13992\ : LocalMux
    port map (
            O => \N__57990\,
            I => comm_data_vld
        );

    \I__13991\ : LocalMux
    port map (
            O => \N__57985\,
            I => comm_data_vld
        );

    \I__13990\ : InMux
    port map (
            O => \N__57970\,
            I => \N__57967\
        );

    \I__13989\ : LocalMux
    port map (
            O => \N__57967\,
            I => \N__57964\
        );

    \I__13988\ : Span4Mux_h
    port map (
            O => \N__57964\,
            I => \N__57961\
        );

    \I__13987\ : Odrv4
    port map (
            O => \N__57961\,
            I => n4_adj_1718
        );

    \I__13986\ : InMux
    port map (
            O => \N__57958\,
            I => \N__57954\
        );

    \I__13985\ : CascadeMux
    port map (
            O => \N__57957\,
            I => \N__57950\
        );

    \I__13984\ : LocalMux
    port map (
            O => \N__57954\,
            I => \N__57947\
        );

    \I__13983\ : InMux
    port map (
            O => \N__57953\,
            I => \N__57942\
        );

    \I__13982\ : InMux
    port map (
            O => \N__57950\,
            I => \N__57942\
        );

    \I__13981\ : Odrv4
    port map (
            O => \N__57947\,
            I => req_data_cnt_11
        );

    \I__13980\ : LocalMux
    port map (
            O => \N__57942\,
            I => req_data_cnt_11
        );

    \I__13979\ : InMux
    port map (
            O => \N__57937\,
            I => \N__57934\
        );

    \I__13978\ : LocalMux
    port map (
            O => \N__57934\,
            I => \N__57931\
        );

    \I__13977\ : Span4Mux_h
    port map (
            O => \N__57931\,
            I => \N__57928\
        );

    \I__13976\ : Span4Mux_h
    port map (
            O => \N__57928\,
            I => \N__57925\
        );

    \I__13975\ : Span4Mux_v
    port map (
            O => \N__57925\,
            I => \N__57922\
        );

    \I__13974\ : Odrv4
    port map (
            O => \N__57922\,
            I => n112_adj_1777
        );

    \I__13973\ : InMux
    port map (
            O => \N__57919\,
            I => \N__57916\
        );

    \I__13972\ : LocalMux
    port map (
            O => \N__57916\,
            I => \N__57913\
        );

    \I__13971\ : Span12Mux_h
    port map (
            O => \N__57913\,
            I => \N__57910\
        );

    \I__13970\ : Odrv12
    port map (
            O => \N__57910\,
            I => \comm_buf_0_7_N_543_5\
        );

    \I__13969\ : InMux
    port map (
            O => \N__57907\,
            I => \N__57900\
        );

    \I__13968\ : InMux
    port map (
            O => \N__57906\,
            I => \N__57900\
        );

    \I__13967\ : InMux
    port map (
            O => \N__57905\,
            I => \N__57897\
        );

    \I__13966\ : LocalMux
    port map (
            O => \N__57900\,
            I => n1373
        );

    \I__13965\ : LocalMux
    port map (
            O => \N__57897\,
            I => n1373
        );

    \I__13964\ : CascadeMux
    port map (
            O => \N__57892\,
            I => \n2_cascade_\
        );

    \I__13963\ : InMux
    port map (
            O => \N__57889\,
            I => \N__57886\
        );

    \I__13962\ : LocalMux
    port map (
            O => \N__57886\,
            I => \N__57883\
        );

    \I__13961\ : Odrv4
    port map (
            O => \N__57883\,
            I => n23342
        );

    \I__13960\ : CascadeMux
    port map (
            O => \N__57880\,
            I => \N__57873\
        );

    \I__13959\ : InMux
    port map (
            O => \N__57879\,
            I => \N__57864\
        );

    \I__13958\ : InMux
    port map (
            O => \N__57878\,
            I => \N__57864\
        );

    \I__13957\ : InMux
    port map (
            O => \N__57877\,
            I => \N__57857\
        );

    \I__13956\ : InMux
    port map (
            O => \N__57876\,
            I => \N__57845\
        );

    \I__13955\ : InMux
    port map (
            O => \N__57873\,
            I => \N__57841\
        );

    \I__13954\ : CascadeMux
    port map (
            O => \N__57872\,
            I => \N__57838\
        );

    \I__13953\ : CascadeMux
    port map (
            O => \N__57871\,
            I => \N__57835\
        );

    \I__13952\ : InMux
    port map (
            O => \N__57870\,
            I => \N__57830\
        );

    \I__13951\ : CascadeMux
    port map (
            O => \N__57869\,
            I => \N__57827\
        );

    \I__13950\ : LocalMux
    port map (
            O => \N__57864\,
            I => \N__57824\
        );

    \I__13949\ : InMux
    port map (
            O => \N__57863\,
            I => \N__57821\
        );

    \I__13948\ : InMux
    port map (
            O => \N__57862\,
            I => \N__57814\
        );

    \I__13947\ : InMux
    port map (
            O => \N__57861\,
            I => \N__57814\
        );

    \I__13946\ : InMux
    port map (
            O => \N__57860\,
            I => \N__57814\
        );

    \I__13945\ : LocalMux
    port map (
            O => \N__57857\,
            I => \N__57811\
        );

    \I__13944\ : InMux
    port map (
            O => \N__57856\,
            I => \N__57808\
        );

    \I__13943\ : CascadeMux
    port map (
            O => \N__57855\,
            I => \N__57805\
        );

    \I__13942\ : CascadeMux
    port map (
            O => \N__57854\,
            I => \N__57802\
        );

    \I__13941\ : InMux
    port map (
            O => \N__57853\,
            I => \N__57799\
        );

    \I__13940\ : InMux
    port map (
            O => \N__57852\,
            I => \N__57794\
        );

    \I__13939\ : InMux
    port map (
            O => \N__57851\,
            I => \N__57794\
        );

    \I__13938\ : InMux
    port map (
            O => \N__57850\,
            I => \N__57789\
        );

    \I__13937\ : InMux
    port map (
            O => \N__57849\,
            I => \N__57789\
        );

    \I__13936\ : InMux
    port map (
            O => \N__57848\,
            I => \N__57786\
        );

    \I__13935\ : LocalMux
    port map (
            O => \N__57845\,
            I => \N__57783\
        );

    \I__13934\ : CascadeMux
    port map (
            O => \N__57844\,
            I => \N__57780\
        );

    \I__13933\ : LocalMux
    port map (
            O => \N__57841\,
            I => \N__57775\
        );

    \I__13932\ : InMux
    port map (
            O => \N__57838\,
            I => \N__57772\
        );

    \I__13931\ : InMux
    port map (
            O => \N__57835\,
            I => \N__57765\
        );

    \I__13930\ : InMux
    port map (
            O => \N__57834\,
            I => \N__57765\
        );

    \I__13929\ : InMux
    port map (
            O => \N__57833\,
            I => \N__57765\
        );

    \I__13928\ : LocalMux
    port map (
            O => \N__57830\,
            I => \N__57760\
        );

    \I__13927\ : InMux
    port map (
            O => \N__57827\,
            I => \N__57757\
        );

    \I__13926\ : Span4Mux_v
    port map (
            O => \N__57824\,
            I => \N__57754\
        );

    \I__13925\ : LocalMux
    port map (
            O => \N__57821\,
            I => \N__57751\
        );

    \I__13924\ : LocalMux
    port map (
            O => \N__57814\,
            I => \N__57748\
        );

    \I__13923\ : Span4Mux_h
    port map (
            O => \N__57811\,
            I => \N__57742\
        );

    \I__13922\ : LocalMux
    port map (
            O => \N__57808\,
            I => \N__57736\
        );

    \I__13921\ : InMux
    port map (
            O => \N__57805\,
            I => \N__57731\
        );

    \I__13920\ : InMux
    port map (
            O => \N__57802\,
            I => \N__57731\
        );

    \I__13919\ : LocalMux
    port map (
            O => \N__57799\,
            I => \N__57723\
        );

    \I__13918\ : LocalMux
    port map (
            O => \N__57794\,
            I => \N__57723\
        );

    \I__13917\ : LocalMux
    port map (
            O => \N__57789\,
            I => \N__57716\
        );

    \I__13916\ : LocalMux
    port map (
            O => \N__57786\,
            I => \N__57716\
        );

    \I__13915\ : Span4Mux_h
    port map (
            O => \N__57783\,
            I => \N__57716\
        );

    \I__13914\ : InMux
    port map (
            O => \N__57780\,
            I => \N__57713\
        );

    \I__13913\ : CascadeMux
    port map (
            O => \N__57779\,
            I => \N__57697\
        );

    \I__13912\ : CascadeMux
    port map (
            O => \N__57778\,
            I => \N__57694\
        );

    \I__13911\ : Span4Mux_h
    port map (
            O => \N__57775\,
            I => \N__57687\
        );

    \I__13910\ : LocalMux
    port map (
            O => \N__57772\,
            I => \N__57687\
        );

    \I__13909\ : LocalMux
    port map (
            O => \N__57765\,
            I => \N__57684\
        );

    \I__13908\ : InMux
    port map (
            O => \N__57764\,
            I => \N__57681\
        );

    \I__13907\ : CascadeMux
    port map (
            O => \N__57763\,
            I => \N__57678\
        );

    \I__13906\ : Span4Mux_v
    port map (
            O => \N__57760\,
            I => \N__57673\
        );

    \I__13905\ : LocalMux
    port map (
            O => \N__57757\,
            I => \N__57673\
        );

    \I__13904\ : Span4Mux_v
    port map (
            O => \N__57754\,
            I => \N__57666\
        );

    \I__13903\ : Span4Mux_v
    port map (
            O => \N__57751\,
            I => \N__57666\
        );

    \I__13902\ : Span4Mux_v
    port map (
            O => \N__57748\,
            I => \N__57666\
        );

    \I__13901\ : CascadeMux
    port map (
            O => \N__57747\,
            I => \N__57662\
        );

    \I__13900\ : CascadeMux
    port map (
            O => \N__57746\,
            I => \N__57658\
        );

    \I__13899\ : InMux
    port map (
            O => \N__57745\,
            I => \N__57655\
        );

    \I__13898\ : Span4Mux_h
    port map (
            O => \N__57742\,
            I => \N__57652\
        );

    \I__13897\ : InMux
    port map (
            O => \N__57741\,
            I => \N__57647\
        );

    \I__13896\ : InMux
    port map (
            O => \N__57740\,
            I => \N__57647\
        );

    \I__13895\ : InMux
    port map (
            O => \N__57739\,
            I => \N__57644\
        );

    \I__13894\ : Span4Mux_h
    port map (
            O => \N__57736\,
            I => \N__57639\
        );

    \I__13893\ : LocalMux
    port map (
            O => \N__57731\,
            I => \N__57639\
        );

    \I__13892\ : InMux
    port map (
            O => \N__57730\,
            I => \N__57632\
        );

    \I__13891\ : InMux
    port map (
            O => \N__57729\,
            I => \N__57632\
        );

    \I__13890\ : InMux
    port map (
            O => \N__57728\,
            I => \N__57632\
        );

    \I__13889\ : Span4Mux_v
    port map (
            O => \N__57723\,
            I => \N__57625\
        );

    \I__13888\ : Span4Mux_v
    port map (
            O => \N__57716\,
            I => \N__57625\
        );

    \I__13887\ : LocalMux
    port map (
            O => \N__57713\,
            I => \N__57625\
        );

    \I__13886\ : InMux
    port map (
            O => \N__57712\,
            I => \N__57622\
        );

    \I__13885\ : CascadeMux
    port map (
            O => \N__57711\,
            I => \N__57614\
        );

    \I__13884\ : CascadeMux
    port map (
            O => \N__57710\,
            I => \N__57611\
        );

    \I__13883\ : CascadeMux
    port map (
            O => \N__57709\,
            I => \N__57607\
        );

    \I__13882\ : CascadeMux
    port map (
            O => \N__57708\,
            I => \N__57604\
        );

    \I__13881\ : CascadeMux
    port map (
            O => \N__57707\,
            I => \N__57600\
        );

    \I__13880\ : InMux
    port map (
            O => \N__57706\,
            I => \N__57591\
        );

    \I__13879\ : InMux
    port map (
            O => \N__57705\,
            I => \N__57591\
        );

    \I__13878\ : InMux
    port map (
            O => \N__57704\,
            I => \N__57591\
        );

    \I__13877\ : InMux
    port map (
            O => \N__57703\,
            I => \N__57591\
        );

    \I__13876\ : InMux
    port map (
            O => \N__57702\,
            I => \N__57588\
        );

    \I__13875\ : CascadeMux
    port map (
            O => \N__57701\,
            I => \N__57584\
        );

    \I__13874\ : InMux
    port map (
            O => \N__57700\,
            I => \N__57571\
        );

    \I__13873\ : InMux
    port map (
            O => \N__57697\,
            I => \N__57571\
        );

    \I__13872\ : InMux
    port map (
            O => \N__57694\,
            I => \N__57571\
        );

    \I__13871\ : InMux
    port map (
            O => \N__57693\,
            I => \N__57571\
        );

    \I__13870\ : InMux
    port map (
            O => \N__57692\,
            I => \N__57571\
        );

    \I__13869\ : Span4Mux_h
    port map (
            O => \N__57687\,
            I => \N__57566\
        );

    \I__13868\ : Span4Mux_h
    port map (
            O => \N__57684\,
            I => \N__57566\
        );

    \I__13867\ : LocalMux
    port map (
            O => \N__57681\,
            I => \N__57563\
        );

    \I__13866\ : InMux
    port map (
            O => \N__57678\,
            I => \N__57560\
        );

    \I__13865\ : Sp12to4
    port map (
            O => \N__57673\,
            I => \N__57557\
        );

    \I__13864\ : Span4Mux_h
    port map (
            O => \N__57666\,
            I => \N__57554\
        );

    \I__13863\ : InMux
    port map (
            O => \N__57665\,
            I => \N__57551\
        );

    \I__13862\ : InMux
    port map (
            O => \N__57662\,
            I => \N__57546\
        );

    \I__13861\ : InMux
    port map (
            O => \N__57661\,
            I => \N__57546\
        );

    \I__13860\ : InMux
    port map (
            O => \N__57658\,
            I => \N__57543\
        );

    \I__13859\ : LocalMux
    port map (
            O => \N__57655\,
            I => \N__57540\
        );

    \I__13858\ : Span4Mux_h
    port map (
            O => \N__57652\,
            I => \N__57535\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__57647\,
            I => \N__57535\
        );

    \I__13856\ : LocalMux
    port map (
            O => \N__57644\,
            I => \N__57532\
        );

    \I__13855\ : Span4Mux_h
    port map (
            O => \N__57639\,
            I => \N__57527\
        );

    \I__13854\ : LocalMux
    port map (
            O => \N__57632\,
            I => \N__57527\
        );

    \I__13853\ : Span4Mux_h
    port map (
            O => \N__57625\,
            I => \N__57522\
        );

    \I__13852\ : LocalMux
    port map (
            O => \N__57622\,
            I => \N__57522\
        );

    \I__13851\ : InMux
    port map (
            O => \N__57621\,
            I => \N__57517\
        );

    \I__13850\ : InMux
    port map (
            O => \N__57620\,
            I => \N__57514\
        );

    \I__13849\ : InMux
    port map (
            O => \N__57619\,
            I => \N__57509\
        );

    \I__13848\ : InMux
    port map (
            O => \N__57618\,
            I => \N__57509\
        );

    \I__13847\ : InMux
    port map (
            O => \N__57617\,
            I => \N__57506\
        );

    \I__13846\ : InMux
    port map (
            O => \N__57614\,
            I => \N__57501\
        );

    \I__13845\ : InMux
    port map (
            O => \N__57611\,
            I => \N__57501\
        );

    \I__13844\ : InMux
    port map (
            O => \N__57610\,
            I => \N__57498\
        );

    \I__13843\ : InMux
    port map (
            O => \N__57607\,
            I => \N__57489\
        );

    \I__13842\ : InMux
    port map (
            O => \N__57604\,
            I => \N__57489\
        );

    \I__13841\ : InMux
    port map (
            O => \N__57603\,
            I => \N__57489\
        );

    \I__13840\ : InMux
    port map (
            O => \N__57600\,
            I => \N__57489\
        );

    \I__13839\ : LocalMux
    port map (
            O => \N__57591\,
            I => \N__57484\
        );

    \I__13838\ : LocalMux
    port map (
            O => \N__57588\,
            I => \N__57484\
        );

    \I__13837\ : InMux
    port map (
            O => \N__57587\,
            I => \N__57475\
        );

    \I__13836\ : InMux
    port map (
            O => \N__57584\,
            I => \N__57475\
        );

    \I__13835\ : InMux
    port map (
            O => \N__57583\,
            I => \N__57475\
        );

    \I__13834\ : InMux
    port map (
            O => \N__57582\,
            I => \N__57475\
        );

    \I__13833\ : LocalMux
    port map (
            O => \N__57571\,
            I => \N__57472\
        );

    \I__13832\ : Sp12to4
    port map (
            O => \N__57566\,
            I => \N__57469\
        );

    \I__13831\ : Span4Mux_h
    port map (
            O => \N__57563\,
            I => \N__57465\
        );

    \I__13830\ : LocalMux
    port map (
            O => \N__57560\,
            I => \N__57462\
        );

    \I__13829\ : Span12Mux_v
    port map (
            O => \N__57557\,
            I => \N__57455\
        );

    \I__13828\ : Sp12to4
    port map (
            O => \N__57554\,
            I => \N__57455\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__57551\,
            I => \N__57455\
        );

    \I__13826\ : LocalMux
    port map (
            O => \N__57546\,
            I => \N__57450\
        );

    \I__13825\ : LocalMux
    port map (
            O => \N__57543\,
            I => \N__57450\
        );

    \I__13824\ : Span4Mux_v
    port map (
            O => \N__57540\,
            I => \N__57445\
        );

    \I__13823\ : Span4Mux_h
    port map (
            O => \N__57535\,
            I => \N__57445\
        );

    \I__13822\ : Span4Mux_h
    port map (
            O => \N__57532\,
            I => \N__57438\
        );

    \I__13821\ : Span4Mux_v
    port map (
            O => \N__57527\,
            I => \N__57438\
        );

    \I__13820\ : Span4Mux_h
    port map (
            O => \N__57522\,
            I => \N__57438\
        );

    \I__13819\ : InMux
    port map (
            O => \N__57521\,
            I => \N__57435\
        );

    \I__13818\ : InMux
    port map (
            O => \N__57520\,
            I => \N__57432\
        );

    \I__13817\ : LocalMux
    port map (
            O => \N__57517\,
            I => \N__57429\
        );

    \I__13816\ : LocalMux
    port map (
            O => \N__57514\,
            I => \N__57408\
        );

    \I__13815\ : LocalMux
    port map (
            O => \N__57509\,
            I => \N__57408\
        );

    \I__13814\ : LocalMux
    port map (
            O => \N__57506\,
            I => \N__57408\
        );

    \I__13813\ : LocalMux
    port map (
            O => \N__57501\,
            I => \N__57408\
        );

    \I__13812\ : LocalMux
    port map (
            O => \N__57498\,
            I => \N__57408\
        );

    \I__13811\ : LocalMux
    port map (
            O => \N__57489\,
            I => \N__57408\
        );

    \I__13810\ : Sp12to4
    port map (
            O => \N__57484\,
            I => \N__57408\
        );

    \I__13809\ : LocalMux
    port map (
            O => \N__57475\,
            I => \N__57408\
        );

    \I__13808\ : Sp12to4
    port map (
            O => \N__57472\,
            I => \N__57408\
        );

    \I__13807\ : Span12Mux_s6_v
    port map (
            O => \N__57469\,
            I => \N__57408\
        );

    \I__13806\ : InMux
    port map (
            O => \N__57468\,
            I => \N__57405\
        );

    \I__13805\ : Span4Mux_h
    port map (
            O => \N__57465\,
            I => \N__57400\
        );

    \I__13804\ : Span4Mux_v
    port map (
            O => \N__57462\,
            I => \N__57400\
        );

    \I__13803\ : Span12Mux_h
    port map (
            O => \N__57455\,
            I => \N__57397\
        );

    \I__13802\ : Span12Mux_h
    port map (
            O => \N__57450\,
            I => \N__57394\
        );

    \I__13801\ : Span4Mux_h
    port map (
            O => \N__57445\,
            I => \N__57389\
        );

    \I__13800\ : Span4Mux_v
    port map (
            O => \N__57438\,
            I => \N__57389\
        );

    \I__13799\ : LocalMux
    port map (
            O => \N__57435\,
            I => \N__57380\
        );

    \I__13798\ : LocalMux
    port map (
            O => \N__57432\,
            I => \N__57380\
        );

    \I__13797\ : Span12Mux_h
    port map (
            O => \N__57429\,
            I => \N__57380\
        );

    \I__13796\ : Span12Mux_v
    port map (
            O => \N__57408\,
            I => \N__57380\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__57405\,
            I => n9837
        );

    \I__13794\ : Odrv4
    port map (
            O => \N__57400\,
            I => n9837
        );

    \I__13793\ : Odrv12
    port map (
            O => \N__57397\,
            I => n9837
        );

    \I__13792\ : Odrv12
    port map (
            O => \N__57394\,
            I => n9837
        );

    \I__13791\ : Odrv4
    port map (
            O => \N__57389\,
            I => n9837
        );

    \I__13790\ : Odrv12
    port map (
            O => \N__57380\,
            I => n9837
        );

    \I__13789\ : CascadeMux
    port map (
            O => \N__57367\,
            I => \n23345_cascade_\
        );

    \I__13788\ : InMux
    port map (
            O => \N__57364\,
            I => \N__57361\
        );

    \I__13787\ : LocalMux
    port map (
            O => \N__57361\,
            I => n8_adj_1659
        );

    \I__13786\ : InMux
    port map (
            O => \N__57358\,
            I => \N__57355\
        );

    \I__13785\ : LocalMux
    port map (
            O => \N__57355\,
            I => \N__57350\
        );

    \I__13784\ : InMux
    port map (
            O => \N__57354\,
            I => \N__57347\
        );

    \I__13783\ : InMux
    port map (
            O => \N__57353\,
            I => \N__57344\
        );

    \I__13782\ : Odrv4
    port map (
            O => \N__57350\,
            I => n2562
        );

    \I__13781\ : LocalMux
    port map (
            O => \N__57347\,
            I => n2562
        );

    \I__13780\ : LocalMux
    port map (
            O => \N__57344\,
            I => n2562
        );

    \I__13779\ : InMux
    port map (
            O => \N__57337\,
            I => \N__57334\
        );

    \I__13778\ : LocalMux
    port map (
            O => \N__57334\,
            I => \N__57331\
        );

    \I__13777\ : Odrv4
    port map (
            O => \N__57331\,
            I => n22339
        );

    \I__13776\ : CascadeMux
    port map (
            O => \N__57328\,
            I => \n22340_cascade_\
        );

    \I__13775\ : CEMux
    port map (
            O => \N__57325\,
            I => \N__57322\
        );

    \I__13774\ : LocalMux
    port map (
            O => \N__57322\,
            I => \N__57319\
        );

    \I__13773\ : Span4Mux_h
    port map (
            O => \N__57319\,
            I => \N__57316\
        );

    \I__13772\ : Span4Mux_h
    port map (
            O => \N__57316\,
            I => \N__57313\
        );

    \I__13771\ : Odrv4
    port map (
            O => \N__57313\,
            I => n14_adj_1593
        );

    \I__13770\ : CascadeMux
    port map (
            O => \N__57310\,
            I => \N__57307\
        );

    \I__13769\ : InMux
    port map (
            O => \N__57307\,
            I => \N__57304\
        );

    \I__13768\ : LocalMux
    port map (
            O => \N__57304\,
            I => \N__57301\
        );

    \I__13767\ : Span4Mux_h
    port map (
            O => \N__57301\,
            I => \N__57296\
        );

    \I__13766\ : InMux
    port map (
            O => \N__57300\,
            I => \N__57293\
        );

    \I__13765\ : InMux
    port map (
            O => \N__57299\,
            I => \N__57290\
        );

    \I__13764\ : Odrv4
    port map (
            O => \N__57296\,
            I => n5
        );

    \I__13763\ : LocalMux
    port map (
            O => \N__57293\,
            I => n5
        );

    \I__13762\ : LocalMux
    port map (
            O => \N__57290\,
            I => n5
        );

    \I__13761\ : CascadeMux
    port map (
            O => \N__57283\,
            I => \n9725_cascade_\
        );

    \I__13760\ : InMux
    port map (
            O => \N__57280\,
            I => \N__57277\
        );

    \I__13759\ : LocalMux
    port map (
            O => \N__57277\,
            I => \N__57274\
        );

    \I__13758\ : Span4Mux_h
    port map (
            O => \N__57274\,
            I => \N__57271\
        );

    \I__13757\ : Odrv4
    port map (
            O => \N__57271\,
            I => n4
        );

    \I__13756\ : InMux
    port map (
            O => \N__57268\,
            I => \N__57265\
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__57265\,
            I => \ADC_VDC.genclk.n28_adj_1481\
        );

    \I__13754\ : CascadeMux
    port map (
            O => \N__57262\,
            I => \N__57258\
        );

    \I__13753\ : InMux
    port map (
            O => \N__57261\,
            I => \N__57255\
        );

    \I__13752\ : InMux
    port map (
            O => \N__57258\,
            I => \N__57252\
        );

    \I__13751\ : LocalMux
    port map (
            O => \N__57255\,
            I => \N__57249\
        );

    \I__13750\ : LocalMux
    port map (
            O => \N__57252\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__13749\ : Odrv4
    port map (
            O => \N__57249\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__13748\ : InMux
    port map (
            O => \N__57244\,
            I => \N__57240\
        );

    \I__13747\ : InMux
    port map (
            O => \N__57243\,
            I => \N__57237\
        );

    \I__13746\ : LocalMux
    port map (
            O => \N__57240\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__13745\ : LocalMux
    port map (
            O => \N__57237\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__13744\ : CascadeMux
    port map (
            O => \N__57232\,
            I => \N__57228\
        );

    \I__13743\ : InMux
    port map (
            O => \N__57231\,
            I => \N__57225\
        );

    \I__13742\ : InMux
    port map (
            O => \N__57228\,
            I => \N__57222\
        );

    \I__13741\ : LocalMux
    port map (
            O => \N__57225\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__13740\ : LocalMux
    port map (
            O => \N__57222\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__13739\ : InMux
    port map (
            O => \N__57217\,
            I => \N__57213\
        );

    \I__13738\ : InMux
    port map (
            O => \N__57216\,
            I => \N__57210\
        );

    \I__13737\ : LocalMux
    port map (
            O => \N__57213\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__13736\ : LocalMux
    port map (
            O => \N__57210\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__13735\ : InMux
    port map (
            O => \N__57205\,
            I => \N__57202\
        );

    \I__13734\ : LocalMux
    port map (
            O => \N__57202\,
            I => \ADC_VDC.genclk.n26_adj_1482\
        );

    \I__13733\ : CEMux
    port map (
            O => \N__57199\,
            I => \N__57196\
        );

    \I__13732\ : LocalMux
    port map (
            O => \N__57196\,
            I => \N__57192\
        );

    \I__13731\ : CEMux
    port map (
            O => \N__57195\,
            I => \N__57189\
        );

    \I__13730\ : Span4Mux_h
    port map (
            O => \N__57192\,
            I => \N__57186\
        );

    \I__13729\ : LocalMux
    port map (
            O => \N__57189\,
            I => \N__57183\
        );

    \I__13728\ : Odrv4
    port map (
            O => \N__57186\,
            I => \ADC_VDC.genclk.div_state_1__N_1480\
        );

    \I__13727\ : Odrv12
    port map (
            O => \N__57183\,
            I => \ADC_VDC.genclk.div_state_1__N_1480\
        );

    \I__13726\ : InMux
    port map (
            O => \N__57178\,
            I => \N__57167\
        );

    \I__13725\ : InMux
    port map (
            O => \N__57177\,
            I => \N__57164\
        );

    \I__13724\ : InMux
    port map (
            O => \N__57176\,
            I => \N__57161\
        );

    \I__13723\ : InMux
    port map (
            O => \N__57175\,
            I => \N__57148\
        );

    \I__13722\ : InMux
    port map (
            O => \N__57174\,
            I => \N__57148\
        );

    \I__13721\ : InMux
    port map (
            O => \N__57173\,
            I => \N__57148\
        );

    \I__13720\ : InMux
    port map (
            O => \N__57172\,
            I => \N__57148\
        );

    \I__13719\ : InMux
    port map (
            O => \N__57171\,
            I => \N__57148\
        );

    \I__13718\ : InMux
    port map (
            O => \N__57170\,
            I => \N__57148\
        );

    \I__13717\ : LocalMux
    port map (
            O => \N__57167\,
            I => \N__57138\
        );

    \I__13716\ : LocalMux
    port map (
            O => \N__57164\,
            I => \N__57138\
        );

    \I__13715\ : LocalMux
    port map (
            O => \N__57161\,
            I => \N__57138\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__57148\,
            I => \N__57138\
        );

    \I__13713\ : CascadeMux
    port map (
            O => \N__57147\,
            I => \N__57132\
        );

    \I__13712\ : Span4Mux_v
    port map (
            O => \N__57138\,
            I => \N__57126\
        );

    \I__13711\ : InMux
    port map (
            O => \N__57137\,
            I => \N__57123\
        );

    \I__13710\ : InMux
    port map (
            O => \N__57136\,
            I => \N__57100\
        );

    \I__13709\ : InMux
    port map (
            O => \N__57135\,
            I => \N__57100\
        );

    \I__13708\ : InMux
    port map (
            O => \N__57132\,
            I => \N__57100\
        );

    \I__13707\ : InMux
    port map (
            O => \N__57131\,
            I => \N__57100\
        );

    \I__13706\ : InMux
    port map (
            O => \N__57130\,
            I => \N__57097\
        );

    \I__13705\ : InMux
    port map (
            O => \N__57129\,
            I => \N__57093\
        );

    \I__13704\ : Span4Mux_h
    port map (
            O => \N__57126\,
            I => \N__57087\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__57123\,
            I => \N__57087\
        );

    \I__13702\ : SRMux
    port map (
            O => \N__57122\,
            I => \N__57084\
        );

    \I__13701\ : InMux
    port map (
            O => \N__57121\,
            I => \N__57079\
        );

    \I__13700\ : InMux
    port map (
            O => \N__57120\,
            I => \N__57079\
        );

    \I__13699\ : InMux
    port map (
            O => \N__57119\,
            I => \N__57074\
        );

    \I__13698\ : InMux
    port map (
            O => \N__57118\,
            I => \N__57071\
        );

    \I__13697\ : InMux
    port map (
            O => \N__57117\,
            I => \N__57063\
        );

    \I__13696\ : InMux
    port map (
            O => \N__57116\,
            I => \N__57063\
        );

    \I__13695\ : InMux
    port map (
            O => \N__57115\,
            I => \N__57063\
        );

    \I__13694\ : InMux
    port map (
            O => \N__57114\,
            I => \N__57058\
        );

    \I__13693\ : InMux
    port map (
            O => \N__57113\,
            I => \N__57058\
        );

    \I__13692\ : InMux
    port map (
            O => \N__57112\,
            I => \N__57053\
        );

    \I__13691\ : InMux
    port map (
            O => \N__57111\,
            I => \N__57053\
        );

    \I__13690\ : InMux
    port map (
            O => \N__57110\,
            I => \N__57050\
        );

    \I__13689\ : InMux
    port map (
            O => \N__57109\,
            I => \N__57046\
        );

    \I__13688\ : LocalMux
    port map (
            O => \N__57100\,
            I => \N__57043\
        );

    \I__13687\ : LocalMux
    port map (
            O => \N__57097\,
            I => \N__57040\
        );

    \I__13686\ : InMux
    port map (
            O => \N__57096\,
            I => \N__57037\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__57093\,
            I => \N__57034\
        );

    \I__13684\ : SRMux
    port map (
            O => \N__57092\,
            I => \N__57031\
        );

    \I__13683\ : Span4Mux_v
    port map (
            O => \N__57087\,
            I => \N__57028\
        );

    \I__13682\ : LocalMux
    port map (
            O => \N__57084\,
            I => \N__57025\
        );

    \I__13681\ : LocalMux
    port map (
            O => \N__57079\,
            I => \N__57022\
        );

    \I__13680\ : SRMux
    port map (
            O => \N__57078\,
            I => \N__57019\
        );

    \I__13679\ : InMux
    port map (
            O => \N__57077\,
            I => \N__57016\
        );

    \I__13678\ : LocalMux
    port map (
            O => \N__57074\,
            I => \N__57011\
        );

    \I__13677\ : LocalMux
    port map (
            O => \N__57071\,
            I => \N__57011\
        );

    \I__13676\ : InMux
    port map (
            O => \N__57070\,
            I => \N__57008\
        );

    \I__13675\ : LocalMux
    port map (
            O => \N__57063\,
            I => \N__57003\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__57058\,
            I => \N__57003\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__57053\,
            I => \N__57000\
        );

    \I__13672\ : LocalMux
    port map (
            O => \N__57050\,
            I => \N__56997\
        );

    \I__13671\ : InMux
    port map (
            O => \N__57049\,
            I => \N__56994\
        );

    \I__13670\ : LocalMux
    port map (
            O => \N__57046\,
            I => \N__56989\
        );

    \I__13669\ : Span4Mux_v
    port map (
            O => \N__57043\,
            I => \N__56989\
        );

    \I__13668\ : Span4Mux_h
    port map (
            O => \N__57040\,
            I => \N__56984\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__57037\,
            I => \N__56984\
        );

    \I__13666\ : Span4Mux_h
    port map (
            O => \N__57034\,
            I => \N__56979\
        );

    \I__13665\ : LocalMux
    port map (
            O => \N__57031\,
            I => \N__56979\
        );

    \I__13664\ : Span4Mux_h
    port map (
            O => \N__57028\,
            I => \N__56972\
        );

    \I__13663\ : Span4Mux_v
    port map (
            O => \N__57025\,
            I => \N__56972\
        );

    \I__13662\ : Span4Mux_v
    port map (
            O => \N__57022\,
            I => \N__56972\
        );

    \I__13661\ : LocalMux
    port map (
            O => \N__57019\,
            I => \N__56969\
        );

    \I__13660\ : LocalMux
    port map (
            O => \N__57016\,
            I => \N__56962\
        );

    \I__13659\ : Span4Mux_v
    port map (
            O => \N__57011\,
            I => \N__56962\
        );

    \I__13658\ : LocalMux
    port map (
            O => \N__57008\,
            I => \N__56962\
        );

    \I__13657\ : Span4Mux_v
    port map (
            O => \N__57003\,
            I => \N__56957\
        );

    \I__13656\ : Span4Mux_v
    port map (
            O => \N__57000\,
            I => \N__56957\
        );

    \I__13655\ : Span4Mux_v
    port map (
            O => \N__56997\,
            I => \N__56950\
        );

    \I__13654\ : LocalMux
    port map (
            O => \N__56994\,
            I => \N__56950\
        );

    \I__13653\ : Span4Mux_h
    port map (
            O => \N__56989\,
            I => \N__56950\
        );

    \I__13652\ : Span4Mux_h
    port map (
            O => \N__56984\,
            I => \N__56947\
        );

    \I__13651\ : Span4Mux_v
    port map (
            O => \N__56979\,
            I => \N__56938\
        );

    \I__13650\ : Span4Mux_h
    port map (
            O => \N__56972\,
            I => \N__56938\
        );

    \I__13649\ : Span4Mux_v
    port map (
            O => \N__56969\,
            I => \N__56938\
        );

    \I__13648\ : Span4Mux_h
    port map (
            O => \N__56962\,
            I => \N__56938\
        );

    \I__13647\ : Span4Mux_h
    port map (
            O => \N__56957\,
            I => \N__56933\
        );

    \I__13646\ : Span4Mux_h
    port map (
            O => \N__56950\,
            I => \N__56933\
        );

    \I__13645\ : Odrv4
    port map (
            O => \N__56947\,
            I => comm_clear
        );

    \I__13644\ : Odrv4
    port map (
            O => \N__56938\,
            I => comm_clear
        );

    \I__13643\ : Odrv4
    port map (
            O => \N__56933\,
            I => comm_clear
        );

    \I__13642\ : InMux
    port map (
            O => \N__56926\,
            I => \N__56923\
        );

    \I__13641\ : LocalMux
    port map (
            O => \N__56923\,
            I => \N__56920\
        );

    \I__13640\ : Odrv4
    port map (
            O => \N__56920\,
            I => buf_data_iac_18
        );

    \I__13639\ : CascadeMux
    port map (
            O => \N__56917\,
            I => \N__56914\
        );

    \I__13638\ : InMux
    port map (
            O => \N__56914\,
            I => \N__56911\
        );

    \I__13637\ : LocalMux
    port map (
            O => \N__56911\,
            I => \N__56908\
        );

    \I__13636\ : Span4Mux_h
    port map (
            O => \N__56908\,
            I => \N__56905\
        );

    \I__13635\ : Span4Mux_h
    port map (
            O => \N__56905\,
            I => \N__56902\
        );

    \I__13634\ : Span4Mux_v
    port map (
            O => \N__56902\,
            I => \N__56899\
        );

    \I__13633\ : Odrv4
    port map (
            O => \N__56899\,
            I => n22170
        );

    \I__13632\ : CEMux
    port map (
            O => \N__56896\,
            I => \N__56893\
        );

    \I__13631\ : LocalMux
    port map (
            O => \N__56893\,
            I => \N__56890\
        );

    \I__13630\ : Span4Mux_h
    port map (
            O => \N__56890\,
            I => \N__56887\
        );

    \I__13629\ : Odrv4
    port map (
            O => \N__56887\,
            I => n12035
        );

    \I__13628\ : InMux
    port map (
            O => \N__56884\,
            I => \N__56881\
        );

    \I__13627\ : LocalMux
    port map (
            O => \N__56881\,
            I => \N__56878\
        );

    \I__13626\ : Odrv12
    port map (
            O => \N__56878\,
            I => n7_adj_1687
        );

    \I__13625\ : InMux
    port map (
            O => \N__56875\,
            I => \N__56872\
        );

    \I__13624\ : LocalMux
    port map (
            O => \N__56872\,
            I => \N__56868\
        );

    \I__13623\ : InMux
    port map (
            O => \N__56871\,
            I => \N__56865\
        );

    \I__13622\ : Span4Mux_h
    port map (
            O => \N__56868\,
            I => \N__56862\
        );

    \I__13621\ : LocalMux
    port map (
            O => \N__56865\,
            I => \N__56859\
        );

    \I__13620\ : Odrv4
    port map (
            O => \N__56862\,
            I => \comm_state_3_N_484_3\
        );

    \I__13619\ : Odrv4
    port map (
            O => \N__56859\,
            I => \comm_state_3_N_484_3\
        );

    \I__13618\ : InMux
    port map (
            O => \N__56854\,
            I => \N__56851\
        );

    \I__13617\ : LocalMux
    port map (
            O => \N__56851\,
            I => \N__56846\
        );

    \I__13616\ : InMux
    port map (
            O => \N__56850\,
            I => \N__56843\
        );

    \I__13615\ : InMux
    port map (
            O => \N__56849\,
            I => \N__56840\
        );

    \I__13614\ : Span4Mux_h
    port map (
            O => \N__56846\,
            I => \N__56835\
        );

    \I__13613\ : LocalMux
    port map (
            O => \N__56843\,
            I => \N__56831\
        );

    \I__13612\ : LocalMux
    port map (
            O => \N__56840\,
            I => \N__56828\
        );

    \I__13611\ : InMux
    port map (
            O => \N__56839\,
            I => \N__56825\
        );

    \I__13610\ : InMux
    port map (
            O => \N__56838\,
            I => \N__56822\
        );

    \I__13609\ : Span4Mux_h
    port map (
            O => \N__56835\,
            I => \N__56819\
        );

    \I__13608\ : InMux
    port map (
            O => \N__56834\,
            I => \N__56816\
        );

    \I__13607\ : Span12Mux_v
    port map (
            O => \N__56831\,
            I => \N__56813\
        );

    \I__13606\ : Span4Mux_h
    port map (
            O => \N__56828\,
            I => \N__56810\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__56825\,
            I => \N__56807\
        );

    \I__13604\ : LocalMux
    port map (
            O => \N__56822\,
            I => \N__56804\
        );

    \I__13603\ : Span4Mux_v
    port map (
            O => \N__56819\,
            I => \N__56799\
        );

    \I__13602\ : LocalMux
    port map (
            O => \N__56816\,
            I => \N__56799\
        );

    \I__13601\ : Span12Mux_h
    port map (
            O => \N__56813\,
            I => \N__56796\
        );

    \I__13600\ : Span4Mux_h
    port map (
            O => \N__56810\,
            I => \N__56793\
        );

    \I__13599\ : Span4Mux_h
    port map (
            O => \N__56807\,
            I => \N__56790\
        );

    \I__13598\ : Span4Mux_v
    port map (
            O => \N__56804\,
            I => \N__56785\
        );

    \I__13597\ : Span4Mux_h
    port map (
            O => \N__56799\,
            I => \N__56785\
        );

    \I__13596\ : Odrv12
    port map (
            O => \N__56796\,
            I => n14_adj_1654
        );

    \I__13595\ : Odrv4
    port map (
            O => \N__56793\,
            I => n14_adj_1654
        );

    \I__13594\ : Odrv4
    port map (
            O => \N__56790\,
            I => n14_adj_1654
        );

    \I__13593\ : Odrv4
    port map (
            O => \N__56785\,
            I => n14_adj_1654
        );

    \I__13592\ : CEMux
    port map (
            O => \N__56776\,
            I => \N__56773\
        );

    \I__13591\ : LocalMux
    port map (
            O => \N__56773\,
            I => \N__56770\
        );

    \I__13590\ : Odrv4
    port map (
            O => \N__56770\,
            I => \ADC_VDC.genclk.n6\
        );

    \I__13589\ : CascadeMux
    port map (
            O => \N__56767\,
            I => \N__56764\
        );

    \I__13588\ : InMux
    port map (
            O => \N__56764\,
            I => \N__56760\
        );

    \I__13587\ : InMux
    port map (
            O => \N__56763\,
            I => \N__56757\
        );

    \I__13586\ : LocalMux
    port map (
            O => \N__56760\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__13585\ : LocalMux
    port map (
            O => \N__56757\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__13584\ : InMux
    port map (
            O => \N__56752\,
            I => \N__56748\
        );

    \I__13583\ : InMux
    port map (
            O => \N__56751\,
            I => \N__56745\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__56748\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__56745\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__13580\ : CascadeMux
    port map (
            O => \N__56740\,
            I => \N__56736\
        );

    \I__13579\ : CascadeMux
    port map (
            O => \N__56739\,
            I => \N__56733\
        );

    \I__13578\ : InMux
    port map (
            O => \N__56736\,
            I => \N__56730\
        );

    \I__13577\ : InMux
    port map (
            O => \N__56733\,
            I => \N__56727\
        );

    \I__13576\ : LocalMux
    port map (
            O => \N__56730\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__13575\ : LocalMux
    port map (
            O => \N__56727\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__13574\ : InMux
    port map (
            O => \N__56722\,
            I => \N__56718\
        );

    \I__13573\ : InMux
    port map (
            O => \N__56721\,
            I => \N__56715\
        );

    \I__13572\ : LocalMux
    port map (
            O => \N__56718\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__13571\ : LocalMux
    port map (
            O => \N__56715\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__13570\ : CascadeMux
    port map (
            O => \N__56710\,
            I => \ADC_VDC.genclk.n22308_cascade_\
        );

    \I__13569\ : InMux
    port map (
            O => \N__56707\,
            I => \N__56703\
        );

    \I__13568\ : InMux
    port map (
            O => \N__56706\,
            I => \N__56700\
        );

    \I__13567\ : LocalMux
    port map (
            O => \N__56703\,
            I => \N__56697\
        );

    \I__13566\ : LocalMux
    port map (
            O => \N__56700\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__13565\ : Odrv4
    port map (
            O => \N__56697\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__13564\ : CascadeMux
    port map (
            O => \N__56692\,
            I => \N__56689\
        );

    \I__13563\ : InMux
    port map (
            O => \N__56689\,
            I => \N__56685\
        );

    \I__13562\ : InMux
    port map (
            O => \N__56688\,
            I => \N__56682\
        );

    \I__13561\ : LocalMux
    port map (
            O => \N__56685\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__13560\ : LocalMux
    port map (
            O => \N__56682\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__13559\ : CascadeMux
    port map (
            O => \N__56677\,
            I => \N__56673\
        );

    \I__13558\ : InMux
    port map (
            O => \N__56676\,
            I => \N__56670\
        );

    \I__13557\ : InMux
    port map (
            O => \N__56673\,
            I => \N__56667\
        );

    \I__13556\ : LocalMux
    port map (
            O => \N__56670\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__13555\ : LocalMux
    port map (
            O => \N__56667\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__13554\ : InMux
    port map (
            O => \N__56662\,
            I => \N__56658\
        );

    \I__13553\ : InMux
    port map (
            O => \N__56661\,
            I => \N__56655\
        );

    \I__13552\ : LocalMux
    port map (
            O => \N__56658\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__13551\ : LocalMux
    port map (
            O => \N__56655\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__13550\ : InMux
    port map (
            O => \N__56650\,
            I => \N__56647\
        );

    \I__13549\ : LocalMux
    port map (
            O => \N__56647\,
            I => \ADC_VDC.genclk.n27_adj_1483\
        );

    \I__13548\ : InMux
    port map (
            O => \N__56644\,
            I => \N__56640\
        );

    \I__13547\ : InMux
    port map (
            O => \N__56643\,
            I => \N__56637\
        );

    \I__13546\ : LocalMux
    port map (
            O => \N__56640\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__13545\ : LocalMux
    port map (
            O => \N__56637\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__13544\ : CascadeMux
    port map (
            O => \N__56632\,
            I => \N__56629\
        );

    \I__13543\ : InMux
    port map (
            O => \N__56629\,
            I => \N__56625\
        );

    \I__13542\ : InMux
    port map (
            O => \N__56628\,
            I => \N__56622\
        );

    \I__13541\ : LocalMux
    port map (
            O => \N__56625\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__13540\ : LocalMux
    port map (
            O => \N__56622\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__13539\ : CascadeMux
    port map (
            O => \N__56617\,
            I => \N__56613\
        );

    \I__13538\ : InMux
    port map (
            O => \N__56616\,
            I => \N__56610\
        );

    \I__13537\ : InMux
    port map (
            O => \N__56613\,
            I => \N__56607\
        );

    \I__13536\ : LocalMux
    port map (
            O => \N__56610\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__13535\ : LocalMux
    port map (
            O => \N__56607\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__13534\ : CascadeMux
    port map (
            O => \N__56602\,
            I => \N__56599\
        );

    \I__13533\ : InMux
    port map (
            O => \N__56599\,
            I => \N__56595\
        );

    \I__13532\ : InMux
    port map (
            O => \N__56598\,
            I => \N__56592\
        );

    \I__13531\ : LocalMux
    port map (
            O => \N__56595\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__13530\ : LocalMux
    port map (
            O => \N__56592\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__13529\ : InMux
    port map (
            O => \N__56587\,
            I => \N__56584\
        );

    \I__13528\ : LocalMux
    port map (
            O => \N__56584\,
            I => \N__56579\
        );

    \I__13527\ : InMux
    port map (
            O => \N__56583\,
            I => \N__56574\
        );

    \I__13526\ : CascadeMux
    port map (
            O => \N__56582\,
            I => \N__56571\
        );

    \I__13525\ : Span4Mux_v
    port map (
            O => \N__56579\,
            I => \N__56566\
        );

    \I__13524\ : InMux
    port map (
            O => \N__56578\,
            I => \N__56563\
        );

    \I__13523\ : InMux
    port map (
            O => \N__56577\,
            I => \N__56560\
        );

    \I__13522\ : LocalMux
    port map (
            O => \N__56574\,
            I => \N__56557\
        );

    \I__13521\ : InMux
    port map (
            O => \N__56571\,
            I => \N__56554\
        );

    \I__13520\ : InMux
    port map (
            O => \N__56570\,
            I => \N__56551\
        );

    \I__13519\ : InMux
    port map (
            O => \N__56569\,
            I => \N__56548\
        );

    \I__13518\ : Span4Mux_h
    port map (
            O => \N__56566\,
            I => \N__56543\
        );

    \I__13517\ : LocalMux
    port map (
            O => \N__56563\,
            I => \N__56543\
        );

    \I__13516\ : LocalMux
    port map (
            O => \N__56560\,
            I => \N__56540\
        );

    \I__13515\ : Span4Mux_v
    port map (
            O => \N__56557\,
            I => \N__56533\
        );

    \I__13514\ : LocalMux
    port map (
            O => \N__56554\,
            I => \N__56533\
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__56551\,
            I => \N__56533\
        );

    \I__13512\ : LocalMux
    port map (
            O => \N__56548\,
            I => \N__56529\
        );

    \I__13511\ : Span4Mux_h
    port map (
            O => \N__56543\,
            I => \N__56526\
        );

    \I__13510\ : Span4Mux_v
    port map (
            O => \N__56540\,
            I => \N__56521\
        );

    \I__13509\ : Span4Mux_h
    port map (
            O => \N__56533\,
            I => \N__56521\
        );

    \I__13508\ : InMux
    port map (
            O => \N__56532\,
            I => \N__56518\
        );

    \I__13507\ : Span12Mux_h
    port map (
            O => \N__56529\,
            I => \N__56515\
        );

    \I__13506\ : Span4Mux_v
    port map (
            O => \N__56526\,
            I => \N__56508\
        );

    \I__13505\ : Span4Mux_h
    port map (
            O => \N__56521\,
            I => \N__56508\
        );

    \I__13504\ : LocalMux
    port map (
            O => \N__56518\,
            I => \N__56508\
        );

    \I__13503\ : Odrv12
    port map (
            O => \N__56515\,
            I => comm_buf_1_5
        );

    \I__13502\ : Odrv4
    port map (
            O => \N__56508\,
            I => comm_buf_1_5
        );

    \I__13501\ : InMux
    port map (
            O => \N__56503\,
            I => \N__56499\
        );

    \I__13500\ : InMux
    port map (
            O => \N__56502\,
            I => \N__56496\
        );

    \I__13499\ : LocalMux
    port map (
            O => \N__56499\,
            I => \N__56490\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__56496\,
            I => \N__56490\
        );

    \I__13497\ : InMux
    port map (
            O => \N__56495\,
            I => \N__56487\
        );

    \I__13496\ : Span12Mux_h
    port map (
            O => \N__56490\,
            I => \N__56484\
        );

    \I__13495\ : LocalMux
    port map (
            O => \N__56487\,
            I => data_index_5
        );

    \I__13494\ : Odrv12
    port map (
            O => \N__56484\,
            I => data_index_5
        );

    \I__13493\ : InMux
    port map (
            O => \N__56479\,
            I => \N__56475\
        );

    \I__13492\ : InMux
    port map (
            O => \N__56478\,
            I => \N__56470\
        );

    \I__13491\ : LocalMux
    port map (
            O => \N__56475\,
            I => \N__56466\
        );

    \I__13490\ : InMux
    port map (
            O => \N__56474\,
            I => \N__56463\
        );

    \I__13489\ : InMux
    port map (
            O => \N__56473\,
            I => \N__56455\
        );

    \I__13488\ : LocalMux
    port map (
            O => \N__56470\,
            I => \N__56452\
        );

    \I__13487\ : InMux
    port map (
            O => \N__56469\,
            I => \N__56448\
        );

    \I__13486\ : Span4Mux_h
    port map (
            O => \N__56466\,
            I => \N__56445\
        );

    \I__13485\ : LocalMux
    port map (
            O => \N__56463\,
            I => \N__56442\
        );

    \I__13484\ : InMux
    port map (
            O => \N__56462\,
            I => \N__56439\
        );

    \I__13483\ : InMux
    port map (
            O => \N__56461\,
            I => \N__56434\
        );

    \I__13482\ : InMux
    port map (
            O => \N__56460\,
            I => \N__56434\
        );

    \I__13481\ : InMux
    port map (
            O => \N__56459\,
            I => \N__56429\
        );

    \I__13480\ : InMux
    port map (
            O => \N__56458\,
            I => \N__56429\
        );

    \I__13479\ : LocalMux
    port map (
            O => \N__56455\,
            I => \N__56426\
        );

    \I__13478\ : Span4Mux_v
    port map (
            O => \N__56452\,
            I => \N__56423\
        );

    \I__13477\ : InMux
    port map (
            O => \N__56451\,
            I => \N__56420\
        );

    \I__13476\ : LocalMux
    port map (
            O => \N__56448\,
            I => \N__56417\
        );

    \I__13475\ : Span4Mux_v
    port map (
            O => \N__56445\,
            I => \N__56414\
        );

    \I__13474\ : Sp12to4
    port map (
            O => \N__56442\,
            I => \N__56405\
        );

    \I__13473\ : LocalMux
    port map (
            O => \N__56439\,
            I => \N__56405\
        );

    \I__13472\ : LocalMux
    port map (
            O => \N__56434\,
            I => \N__56405\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__56429\,
            I => \N__56405\
        );

    \I__13470\ : Span4Mux_v
    port map (
            O => \N__56426\,
            I => \N__56396\
        );

    \I__13469\ : Span4Mux_h
    port map (
            O => \N__56423\,
            I => \N__56396\
        );

    \I__13468\ : LocalMux
    port map (
            O => \N__56420\,
            I => \N__56396\
        );

    \I__13467\ : Span4Mux_h
    port map (
            O => \N__56417\,
            I => \N__56396\
        );

    \I__13466\ : Odrv4
    port map (
            O => \N__56414\,
            I => n9324
        );

    \I__13465\ : Odrv12
    port map (
            O => \N__56405\,
            I => n9324
        );

    \I__13464\ : Odrv4
    port map (
            O => \N__56396\,
            I => n9324
        );

    \I__13463\ : InMux
    port map (
            O => \N__56389\,
            I => \N__56386\
        );

    \I__13462\ : LocalMux
    port map (
            O => \N__56386\,
            I => n8_adj_1623
        );

    \I__13461\ : CascadeMux
    port map (
            O => \N__56383\,
            I => \n8_adj_1623_cascade_\
        );

    \I__13460\ : CascadeMux
    port map (
            O => \N__56380\,
            I => \N__56377\
        );

    \I__13459\ : InMux
    port map (
            O => \N__56377\,
            I => \N__56373\
        );

    \I__13458\ : InMux
    port map (
            O => \N__56376\,
            I => \N__56370\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__56373\,
            I => \N__56365\
        );

    \I__13456\ : LocalMux
    port map (
            O => \N__56370\,
            I => \N__56365\
        );

    \I__13455\ : Odrv12
    port map (
            O => \N__56365\,
            I => n7_adj_1622
        );

    \I__13454\ : CascadeMux
    port map (
            O => \N__56362\,
            I => \N__56359\
        );

    \I__13453\ : CascadeBuf
    port map (
            O => \N__56359\,
            I => \N__56356\
        );

    \I__13452\ : CascadeMux
    port map (
            O => \N__56356\,
            I => \N__56353\
        );

    \I__13451\ : CascadeBuf
    port map (
            O => \N__56353\,
            I => \N__56350\
        );

    \I__13450\ : CascadeMux
    port map (
            O => \N__56350\,
            I => \N__56347\
        );

    \I__13449\ : CascadeBuf
    port map (
            O => \N__56347\,
            I => \N__56344\
        );

    \I__13448\ : CascadeMux
    port map (
            O => \N__56344\,
            I => \N__56341\
        );

    \I__13447\ : CascadeBuf
    port map (
            O => \N__56341\,
            I => \N__56338\
        );

    \I__13446\ : CascadeMux
    port map (
            O => \N__56338\,
            I => \N__56335\
        );

    \I__13445\ : CascadeBuf
    port map (
            O => \N__56335\,
            I => \N__56332\
        );

    \I__13444\ : CascadeMux
    port map (
            O => \N__56332\,
            I => \N__56329\
        );

    \I__13443\ : CascadeBuf
    port map (
            O => \N__56329\,
            I => \N__56325\
        );

    \I__13442\ : CascadeMux
    port map (
            O => \N__56328\,
            I => \N__56322\
        );

    \I__13441\ : CascadeMux
    port map (
            O => \N__56325\,
            I => \N__56319\
        );

    \I__13440\ : CascadeBuf
    port map (
            O => \N__56322\,
            I => \N__56316\
        );

    \I__13439\ : CascadeBuf
    port map (
            O => \N__56319\,
            I => \N__56313\
        );

    \I__13438\ : CascadeMux
    port map (
            O => \N__56316\,
            I => \N__56310\
        );

    \I__13437\ : CascadeMux
    port map (
            O => \N__56313\,
            I => \N__56307\
        );

    \I__13436\ : InMux
    port map (
            O => \N__56310\,
            I => \N__56304\
        );

    \I__13435\ : CascadeBuf
    port map (
            O => \N__56307\,
            I => \N__56301\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__56304\,
            I => \N__56298\
        );

    \I__13433\ : CascadeMux
    port map (
            O => \N__56301\,
            I => \N__56295\
        );

    \I__13432\ : Span4Mux_h
    port map (
            O => \N__56298\,
            I => \N__56292\
        );

    \I__13431\ : CascadeBuf
    port map (
            O => \N__56295\,
            I => \N__56289\
        );

    \I__13430\ : Span4Mux_v
    port map (
            O => \N__56292\,
            I => \N__56286\
        );

    \I__13429\ : CascadeMux
    port map (
            O => \N__56289\,
            I => \N__56283\
        );

    \I__13428\ : Span4Mux_v
    port map (
            O => \N__56286\,
            I => \N__56280\
        );

    \I__13427\ : InMux
    port map (
            O => \N__56283\,
            I => \N__56277\
        );

    \I__13426\ : Span4Mux_h
    port map (
            O => \N__56280\,
            I => \N__56274\
        );

    \I__13425\ : LocalMux
    port map (
            O => \N__56277\,
            I => \N__56271\
        );

    \I__13424\ : Span4Mux_h
    port map (
            O => \N__56274\,
            I => \N__56268\
        );

    \I__13423\ : Span4Mux_h
    port map (
            O => \N__56271\,
            I => \N__56265\
        );

    \I__13422\ : Span4Mux_h
    port map (
            O => \N__56268\,
            I => \N__56260\
        );

    \I__13421\ : Span4Mux_v
    port map (
            O => \N__56265\,
            I => \N__56260\
        );

    \I__13420\ : Odrv4
    port map (
            O => \N__56260\,
            I => \data_index_9_N_236_5\
        );

    \I__13419\ : InMux
    port map (
            O => \N__56257\,
            I => \N__56254\
        );

    \I__13418\ : LocalMux
    port map (
            O => \N__56254\,
            I => \N__56251\
        );

    \I__13417\ : Span4Mux_h
    port map (
            O => \N__56251\,
            I => \N__56248\
        );

    \I__13416\ : Span4Mux_v
    port map (
            O => \N__56248\,
            I => \N__56244\
        );

    \I__13415\ : InMux
    port map (
            O => \N__56247\,
            I => \N__56241\
        );

    \I__13414\ : Odrv4
    port map (
            O => \N__56244\,
            I => n21966
        );

    \I__13413\ : LocalMux
    port map (
            O => \N__56241\,
            I => n21966
        );

    \I__13412\ : CascadeMux
    port map (
            O => \N__56236\,
            I => \N__56233\
        );

    \I__13411\ : InMux
    port map (
            O => \N__56233\,
            I => \N__56229\
        );

    \I__13410\ : CascadeMux
    port map (
            O => \N__56232\,
            I => \N__56225\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__56229\,
            I => \N__56222\
        );

    \I__13408\ : InMux
    port map (
            O => \N__56228\,
            I => \N__56217\
        );

    \I__13407\ : InMux
    port map (
            O => \N__56225\,
            I => \N__56217\
        );

    \I__13406\ : Span4Mux_v
    port map (
            O => \N__56222\,
            I => \N__56212\
        );

    \I__13405\ : LocalMux
    port map (
            O => \N__56217\,
            I => \N__56212\
        );

    \I__13404\ : Span4Mux_v
    port map (
            O => \N__56212\,
            I => \N__56209\
        );

    \I__13403\ : Span4Mux_h
    port map (
            O => \N__56209\,
            I => \N__56206\
        );

    \I__13402\ : Sp12to4
    port map (
            O => \N__56206\,
            I => \N__56202\
        );

    \I__13401\ : CascadeMux
    port map (
            O => \N__56205\,
            I => \N__56199\
        );

    \I__13400\ : Span12Mux_h
    port map (
            O => \N__56202\,
            I => \N__56196\
        );

    \I__13399\ : InMux
    port map (
            O => \N__56199\,
            I => \N__56193\
        );

    \I__13398\ : Span12Mux_v
    port map (
            O => \N__56196\,
            I => \N__56190\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__56193\,
            I => trig_dds1
        );

    \I__13396\ : Odrv12
    port map (
            O => \N__56190\,
            I => trig_dds1
        );

    \I__13395\ : InMux
    port map (
            O => \N__56185\,
            I => \N__56181\
        );

    \I__13394\ : InMux
    port map (
            O => \N__56184\,
            I => \N__56178\
        );

    \I__13393\ : LocalMux
    port map (
            O => \N__56181\,
            I => n21920
        );

    \I__13392\ : LocalMux
    port map (
            O => \N__56178\,
            I => n21920
        );

    \I__13391\ : CascadeMux
    port map (
            O => \N__56173\,
            I => \n22399_cascade_\
        );

    \I__13390\ : InMux
    port map (
            O => \N__56170\,
            I => \N__56167\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__56167\,
            I => \N__56164\
        );

    \I__13388\ : Span4Mux_h
    port map (
            O => \N__56164\,
            I => \N__56161\
        );

    \I__13387\ : Odrv4
    port map (
            O => \N__56161\,
            I => n40_adj_1689
        );

    \I__13386\ : InMux
    port map (
            O => \N__56158\,
            I => \N__56154\
        );

    \I__13385\ : CascadeMux
    port map (
            O => \N__56157\,
            I => \N__56151\
        );

    \I__13384\ : LocalMux
    port map (
            O => \N__56154\,
            I => \N__56148\
        );

    \I__13383\ : InMux
    port map (
            O => \N__56151\,
            I => \N__56145\
        );

    \I__13382\ : Span4Mux_h
    port map (
            O => \N__56148\,
            I => \N__56142\
        );

    \I__13381\ : LocalMux
    port map (
            O => \N__56145\,
            I => data_idxvec_11
        );

    \I__13380\ : Odrv4
    port map (
            O => \N__56142\,
            I => data_idxvec_11
        );

    \I__13379\ : InMux
    port map (
            O => \N__56137\,
            I => \N__56134\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__56134\,
            I => \N__56129\
        );

    \I__13377\ : InMux
    port map (
            O => \N__56133\,
            I => \N__56126\
        );

    \I__13376\ : InMux
    port map (
            O => \N__56132\,
            I => \N__56123\
        );

    \I__13375\ : Span4Mux_v
    port map (
            O => \N__56129\,
            I => \N__56120\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__56126\,
            I => \N__56117\
        );

    \I__13373\ : LocalMux
    port map (
            O => \N__56123\,
            I => data_cntvec_11
        );

    \I__13372\ : Odrv4
    port map (
            O => \N__56120\,
            I => data_cntvec_11
        );

    \I__13371\ : Odrv4
    port map (
            O => \N__56117\,
            I => data_cntvec_11
        );

    \I__13370\ : InMux
    port map (
            O => \N__56110\,
            I => \N__56106\
        );

    \I__13369\ : CascadeMux
    port map (
            O => \N__56109\,
            I => \N__56103\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__56106\,
            I => \N__56100\
        );

    \I__13367\ : InMux
    port map (
            O => \N__56103\,
            I => \N__56097\
        );

    \I__13366\ : Span4Mux_v
    port map (
            O => \N__56100\,
            I => \N__56093\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__56097\,
            I => \N__56090\
        );

    \I__13364\ : InMux
    port map (
            O => \N__56096\,
            I => \N__56087\
        );

    \I__13363\ : Span4Mux_h
    port map (
            O => \N__56093\,
            I => \N__56079\
        );

    \I__13362\ : Span4Mux_v
    port map (
            O => \N__56090\,
            I => \N__56079\
        );

    \I__13361\ : LocalMux
    port map (
            O => \N__56087\,
            I => \N__56079\
        );

    \I__13360\ : CascadeMux
    port map (
            O => \N__56086\,
            I => \N__56075\
        );

    \I__13359\ : Span4Mux_h
    port map (
            O => \N__56079\,
            I => \N__56071\
        );

    \I__13358\ : CascadeMux
    port map (
            O => \N__56078\,
            I => \N__56066\
        );

    \I__13357\ : InMux
    port map (
            O => \N__56075\,
            I => \N__56062\
        );

    \I__13356\ : InMux
    port map (
            O => \N__56074\,
            I => \N__56059\
        );

    \I__13355\ : Span4Mux_h
    port map (
            O => \N__56071\,
            I => \N__56056\
        );

    \I__13354\ : InMux
    port map (
            O => \N__56070\,
            I => \N__56051\
        );

    \I__13353\ : InMux
    port map (
            O => \N__56069\,
            I => \N__56051\
        );

    \I__13352\ : InMux
    port map (
            O => \N__56066\,
            I => \N__56048\
        );

    \I__13351\ : InMux
    port map (
            O => \N__56065\,
            I => \N__56045\
        );

    \I__13350\ : LocalMux
    port map (
            O => \N__56062\,
            I => \N__56042\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__56059\,
            I => \N__56037\
        );

    \I__13348\ : Span4Mux_v
    port map (
            O => \N__56056\,
            I => \N__56037\
        );

    \I__13347\ : LocalMux
    port map (
            O => \N__56051\,
            I => \N__56030\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__56048\,
            I => \N__56030\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__56045\,
            I => \N__56030\
        );

    \I__13344\ : Odrv4
    port map (
            O => \N__56042\,
            I => comm_buf_1_4
        );

    \I__13343\ : Odrv4
    port map (
            O => \N__56037\,
            I => comm_buf_1_4
        );

    \I__13342\ : Odrv12
    port map (
            O => \N__56030\,
            I => comm_buf_1_4
        );

    \I__13341\ : InMux
    port map (
            O => \N__56023\,
            I => \N__56019\
        );

    \I__13340\ : InMux
    port map (
            O => \N__56022\,
            I => \N__56016\
        );

    \I__13339\ : LocalMux
    port map (
            O => \N__56019\,
            I => \N__56013\
        );

    \I__13338\ : LocalMux
    port map (
            O => \N__56016\,
            I => \N__56010\
        );

    \I__13337\ : Span4Mux_h
    port map (
            O => \N__56013\,
            I => \N__56007\
        );

    \I__13336\ : Span4Mux_h
    port map (
            O => \N__56010\,
            I => \N__56004\
        );

    \I__13335\ : Odrv4
    port map (
            O => \N__56007\,
            I => n14_adj_1611
        );

    \I__13334\ : Odrv4
    port map (
            O => \N__56004\,
            I => n14_adj_1611
        );

    \I__13333\ : InMux
    port map (
            O => \N__55999\,
            I => \N__55996\
        );

    \I__13332\ : LocalMux
    port map (
            O => \N__55996\,
            I => \N__55993\
        );

    \I__13331\ : Span4Mux_v
    port map (
            O => \N__55993\,
            I => \N__55990\
        );

    \I__13330\ : Sp12to4
    port map (
            O => \N__55990\,
            I => \N__55987\
        );

    \I__13329\ : Span12Mux_h
    port map (
            O => \N__55987\,
            I => \N__55984\
        );

    \I__13328\ : Odrv12
    port map (
            O => \N__55984\,
            I => n22272
        );

    \I__13327\ : CascadeMux
    port map (
            O => \N__55981\,
            I => \n23420_cascade_\
        );

    \I__13326\ : InMux
    port map (
            O => \N__55978\,
            I => \N__55975\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__55975\,
            I => \N__55972\
        );

    \I__13324\ : Span4Mux_h
    port map (
            O => \N__55972\,
            I => \N__55969\
        );

    \I__13323\ : Odrv4
    port map (
            O => \N__55969\,
            I => n22271
        );

    \I__13322\ : InMux
    port map (
            O => \N__55966\,
            I => \N__55963\
        );

    \I__13321\ : LocalMux
    port map (
            O => \N__55963\,
            I => \N__55960\
        );

    \I__13320\ : Span4Mux_v
    port map (
            O => \N__55960\,
            I => \N__55957\
        );

    \I__13319\ : Span4Mux_v
    port map (
            O => \N__55957\,
            I => \N__55954\
        );

    \I__13318\ : Sp12to4
    port map (
            O => \N__55954\,
            I => \N__55951\
        );

    \I__13317\ : Odrv12
    port map (
            O => \N__55951\,
            I => n111_adj_1719
        );

    \I__13316\ : CascadeMux
    port map (
            O => \N__55948\,
            I => \n23423_cascade_\
        );

    \I__13315\ : CascadeMux
    port map (
            O => \N__55945\,
            I => \N__55942\
        );

    \I__13314\ : InMux
    port map (
            O => \N__55942\,
            I => \N__55938\
        );

    \I__13313\ : CascadeMux
    port map (
            O => \N__55941\,
            I => \N__55932\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__55938\,
            I => \N__55928\
        );

    \I__13311\ : InMux
    port map (
            O => \N__55937\,
            I => \N__55925\
        );

    \I__13310\ : CascadeMux
    port map (
            O => \N__55936\,
            I => \N__55922\
        );

    \I__13309\ : InMux
    port map (
            O => \N__55935\,
            I => \N__55917\
        );

    \I__13308\ : InMux
    port map (
            O => \N__55932\,
            I => \N__55917\
        );

    \I__13307\ : CascadeMux
    port map (
            O => \N__55931\,
            I => \N__55914\
        );

    \I__13306\ : Span4Mux_v
    port map (
            O => \N__55928\,
            I => \N__55909\
        );

    \I__13305\ : LocalMux
    port map (
            O => \N__55925\,
            I => \N__55909\
        );

    \I__13304\ : InMux
    port map (
            O => \N__55922\,
            I => \N__55906\
        );

    \I__13303\ : LocalMux
    port map (
            O => \N__55917\,
            I => \N__55903\
        );

    \I__13302\ : InMux
    port map (
            O => \N__55914\,
            I => \N__55900\
        );

    \I__13301\ : Span4Mux_v
    port map (
            O => \N__55909\,
            I => \N__55896\
        );

    \I__13300\ : LocalMux
    port map (
            O => \N__55906\,
            I => \N__55893\
        );

    \I__13299\ : Span4Mux_v
    port map (
            O => \N__55903\,
            I => \N__55888\
        );

    \I__13298\ : LocalMux
    port map (
            O => \N__55900\,
            I => \N__55888\
        );

    \I__13297\ : InMux
    port map (
            O => \N__55899\,
            I => \N__55885\
        );

    \I__13296\ : Span4Mux_h
    port map (
            O => \N__55896\,
            I => \N__55881\
        );

    \I__13295\ : Span4Mux_v
    port map (
            O => \N__55893\,
            I => \N__55878\
        );

    \I__13294\ : Span4Mux_h
    port map (
            O => \N__55888\,
            I => \N__55873\
        );

    \I__13293\ : LocalMux
    port map (
            O => \N__55885\,
            I => \N__55873\
        );

    \I__13292\ : InMux
    port map (
            O => \N__55884\,
            I => \N__55870\
        );

    \I__13291\ : Span4Mux_h
    port map (
            O => \N__55881\,
            I => \N__55867\
        );

    \I__13290\ : Span4Mux_h
    port map (
            O => \N__55878\,
            I => \N__55862\
        );

    \I__13289\ : Span4Mux_v
    port map (
            O => \N__55873\,
            I => \N__55862\
        );

    \I__13288\ : LocalMux
    port map (
            O => \N__55870\,
            I => \N__55859\
        );

    \I__13287\ : Odrv4
    port map (
            O => \N__55867\,
            I => comm_rx_buf_7
        );

    \I__13286\ : Odrv4
    port map (
            O => \N__55862\,
            I => comm_rx_buf_7
        );

    \I__13285\ : Odrv4
    port map (
            O => \N__55859\,
            I => comm_rx_buf_7
        );

    \I__13284\ : CascadeMux
    port map (
            O => \N__55852\,
            I => \comm_buf_1_7_N_559_7_cascade_\
        );

    \I__13283\ : CascadeMux
    port map (
            O => \N__55849\,
            I => \N__55845\
        );

    \I__13282\ : InMux
    port map (
            O => \N__55848\,
            I => \N__55842\
        );

    \I__13281\ : InMux
    port map (
            O => \N__55845\,
            I => \N__55838\
        );

    \I__13280\ : LocalMux
    port map (
            O => \N__55842\,
            I => \N__55834\
        );

    \I__13279\ : InMux
    port map (
            O => \N__55841\,
            I => \N__55831\
        );

    \I__13278\ : LocalMux
    port map (
            O => \N__55838\,
            I => \N__55828\
        );

    \I__13277\ : CascadeMux
    port map (
            O => \N__55837\,
            I => \N__55824\
        );

    \I__13276\ : Span4Mux_v
    port map (
            O => \N__55834\,
            I => \N__55817\
        );

    \I__13275\ : LocalMux
    port map (
            O => \N__55831\,
            I => \N__55817\
        );

    \I__13274\ : Sp12to4
    port map (
            O => \N__55828\,
            I => \N__55814\
        );

    \I__13273\ : InMux
    port map (
            O => \N__55827\,
            I => \N__55811\
        );

    \I__13272\ : InMux
    port map (
            O => \N__55824\,
            I => \N__55808\
        );

    \I__13271\ : InMux
    port map (
            O => \N__55823\,
            I => \N__55805\
        );

    \I__13270\ : InMux
    port map (
            O => \N__55822\,
            I => \N__55802\
        );

    \I__13269\ : Span4Mux_h
    port map (
            O => \N__55817\,
            I => \N__55799\
        );

    \I__13268\ : Span12Mux_v
    port map (
            O => \N__55814\,
            I => \N__55792\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__55811\,
            I => \N__55792\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__55808\,
            I => \N__55792\
        );

    \I__13265\ : LocalMux
    port map (
            O => \N__55805\,
            I => \N__55787\
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__55802\,
            I => \N__55787\
        );

    \I__13263\ : Span4Mux_h
    port map (
            O => \N__55799\,
            I => \N__55784\
        );

    \I__13262\ : Span12Mux_h
    port map (
            O => \N__55792\,
            I => \N__55781\
        );

    \I__13261\ : Odrv12
    port map (
            O => \N__55787\,
            I => comm_buf_1_7
        );

    \I__13260\ : Odrv4
    port map (
            O => \N__55784\,
            I => comm_buf_1_7
        );

    \I__13259\ : Odrv12
    port map (
            O => \N__55781\,
            I => comm_buf_1_7
        );

    \I__13258\ : CEMux
    port map (
            O => \N__55774\,
            I => \N__55771\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__55771\,
            I => \N__55764\
        );

    \I__13256\ : CEMux
    port map (
            O => \N__55770\,
            I => \N__55761\
        );

    \I__13255\ : CEMux
    port map (
            O => \N__55769\,
            I => \N__55758\
        );

    \I__13254\ : CEMux
    port map (
            O => \N__55768\,
            I => \N__55755\
        );

    \I__13253\ : CEMux
    port map (
            O => \N__55767\,
            I => \N__55752\
        );

    \I__13252\ : Span4Mux_v
    port map (
            O => \N__55764\,
            I => \N__55746\
        );

    \I__13251\ : LocalMux
    port map (
            O => \N__55761\,
            I => \N__55746\
        );

    \I__13250\ : LocalMux
    port map (
            O => \N__55758\,
            I => \N__55743\
        );

    \I__13249\ : LocalMux
    port map (
            O => \N__55755\,
            I => \N__55740\
        );

    \I__13248\ : LocalMux
    port map (
            O => \N__55752\,
            I => \N__55737\
        );

    \I__13247\ : CEMux
    port map (
            O => \N__55751\,
            I => \N__55734\
        );

    \I__13246\ : Span4Mux_h
    port map (
            O => \N__55746\,
            I => \N__55729\
        );

    \I__13245\ : Span4Mux_h
    port map (
            O => \N__55743\,
            I => \N__55729\
        );

    \I__13244\ : Span4Mux_v
    port map (
            O => \N__55740\,
            I => \N__55724\
        );

    \I__13243\ : Span4Mux_h
    port map (
            O => \N__55737\,
            I => \N__55724\
        );

    \I__13242\ : LocalMux
    port map (
            O => \N__55734\,
            I => \N__55721\
        );

    \I__13241\ : Odrv4
    port map (
            O => \N__55729\,
            I => n12761
        );

    \I__13240\ : Odrv4
    port map (
            O => \N__55724\,
            I => n12761
        );

    \I__13239\ : Odrv12
    port map (
            O => \N__55721\,
            I => n12761
        );

    \I__13238\ : SRMux
    port map (
            O => \N__55714\,
            I => \N__55711\
        );

    \I__13237\ : LocalMux
    port map (
            O => \N__55711\,
            I => \N__55704\
        );

    \I__13236\ : SRMux
    port map (
            O => \N__55710\,
            I => \N__55701\
        );

    \I__13235\ : SRMux
    port map (
            O => \N__55709\,
            I => \N__55697\
        );

    \I__13234\ : SRMux
    port map (
            O => \N__55708\,
            I => \N__55694\
        );

    \I__13233\ : SRMux
    port map (
            O => \N__55707\,
            I => \N__55691\
        );

    \I__13232\ : Span4Mux_h
    port map (
            O => \N__55704\,
            I => \N__55686\
        );

    \I__13231\ : LocalMux
    port map (
            O => \N__55701\,
            I => \N__55686\
        );

    \I__13230\ : SRMux
    port map (
            O => \N__55700\,
            I => \N__55683\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__55697\,
            I => \N__55678\
        );

    \I__13228\ : LocalMux
    port map (
            O => \N__55694\,
            I => \N__55678\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__55691\,
            I => \N__55675\
        );

    \I__13226\ : Span4Mux_h
    port map (
            O => \N__55686\,
            I => \N__55670\
        );

    \I__13225\ : LocalMux
    port map (
            O => \N__55683\,
            I => \N__55670\
        );

    \I__13224\ : Span4Mux_v
    port map (
            O => \N__55678\,
            I => \N__55667\
        );

    \I__13223\ : Span4Mux_h
    port map (
            O => \N__55675\,
            I => \N__55664\
        );

    \I__13222\ : Span4Mux_v
    port map (
            O => \N__55670\,
            I => \N__55661\
        );

    \I__13221\ : Span4Mux_h
    port map (
            O => \N__55667\,
            I => \N__55658\
        );

    \I__13220\ : Odrv4
    port map (
            O => \N__55664\,
            I => n15489
        );

    \I__13219\ : Odrv4
    port map (
            O => \N__55661\,
            I => n15489
        );

    \I__13218\ : Odrv4
    port map (
            O => \N__55658\,
            I => n15489
        );

    \I__13217\ : CascadeMux
    port map (
            O => \N__55651\,
            I => \N__55646\
        );

    \I__13216\ : InMux
    port map (
            O => \N__55650\,
            I => \N__55641\
        );

    \I__13215\ : InMux
    port map (
            O => \N__55649\,
            I => \N__55641\
        );

    \I__13214\ : InMux
    port map (
            O => \N__55646\,
            I => \N__55637\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__55641\,
            I => \N__55631\
        );

    \I__13212\ : InMux
    port map (
            O => \N__55640\,
            I => \N__55627\
        );

    \I__13211\ : LocalMux
    port map (
            O => \N__55637\,
            I => \N__55623\
        );

    \I__13210\ : InMux
    port map (
            O => \N__55636\,
            I => \N__55616\
        );

    \I__13209\ : InMux
    port map (
            O => \N__55635\,
            I => \N__55616\
        );

    \I__13208\ : InMux
    port map (
            O => \N__55634\,
            I => \N__55616\
        );

    \I__13207\ : Span4Mux_h
    port map (
            O => \N__55631\,
            I => \N__55613\
        );

    \I__13206\ : InMux
    port map (
            O => \N__55630\,
            I => \N__55610\
        );

    \I__13205\ : LocalMux
    port map (
            O => \N__55627\,
            I => \N__55607\
        );

    \I__13204\ : InMux
    port map (
            O => \N__55626\,
            I => \N__55604\
        );

    \I__13203\ : Span4Mux_v
    port map (
            O => \N__55623\,
            I => \N__55599\
        );

    \I__13202\ : LocalMux
    port map (
            O => \N__55616\,
            I => \N__55599\
        );

    \I__13201\ : Span4Mux_h
    port map (
            O => \N__55613\,
            I => \N__55595\
        );

    \I__13200\ : LocalMux
    port map (
            O => \N__55610\,
            I => \N__55592\
        );

    \I__13199\ : Span4Mux_h
    port map (
            O => \N__55607\,
            I => \N__55589\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__55604\,
            I => \N__55584\
        );

    \I__13197\ : Sp12to4
    port map (
            O => \N__55599\,
            I => \N__55584\
        );

    \I__13196\ : InMux
    port map (
            O => \N__55598\,
            I => \N__55581\
        );

    \I__13195\ : Span4Mux_v
    port map (
            O => \N__55595\,
            I => \N__55576\
        );

    \I__13194\ : Span4Mux_v
    port map (
            O => \N__55592\,
            I => \N__55576\
        );

    \I__13193\ : Span4Mux_v
    port map (
            O => \N__55589\,
            I => \N__55573\
        );

    \I__13192\ : Span12Mux_v
    port map (
            O => \N__55584\,
            I => \N__55570\
        );

    \I__13191\ : LocalMux
    port map (
            O => \N__55581\,
            I => \N__55565\
        );

    \I__13190\ : Span4Mux_h
    port map (
            O => \N__55576\,
            I => \N__55565\
        );

    \I__13189\ : Odrv4
    port map (
            O => \N__55573\,
            I => n18955
        );

    \I__13188\ : Odrv12
    port map (
            O => \N__55570\,
            I => n18955
        );

    \I__13187\ : Odrv4
    port map (
            O => \N__55565\,
            I => n18955
        );

    \I__13186\ : InMux
    port map (
            O => \N__55558\,
            I => \N__55555\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__55555\,
            I => \N__55552\
        );

    \I__13184\ : Odrv4
    port map (
            O => \N__55552\,
            I => n22356
        );

    \I__13183\ : InMux
    port map (
            O => \N__55549\,
            I => \N__55545\
        );

    \I__13182\ : CascadeMux
    port map (
            O => \N__55548\,
            I => \N__55542\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__55545\,
            I => \N__55539\
        );

    \I__13180\ : InMux
    port map (
            O => \N__55542\,
            I => \N__55536\
        );

    \I__13179\ : Span4Mux_v
    port map (
            O => \N__55539\,
            I => \N__55533\
        );

    \I__13178\ : LocalMux
    port map (
            O => \N__55536\,
            I => \N__55530\
        );

    \I__13177\ : Span4Mux_h
    port map (
            O => \N__55533\,
            I => \N__55526\
        );

    \I__13176\ : Span4Mux_v
    port map (
            O => \N__55530\,
            I => \N__55523\
        );

    \I__13175\ : InMux
    port map (
            O => \N__55529\,
            I => \N__55520\
        );

    \I__13174\ : Span4Mux_v
    port map (
            O => \N__55526\,
            I => \N__55515\
        );

    \I__13173\ : Span4Mux_h
    port map (
            O => \N__55523\,
            I => \N__55515\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__55520\,
            I => buf_dds0_13
        );

    \I__13171\ : Odrv4
    port map (
            O => \N__55515\,
            I => buf_dds0_13
        );

    \I__13170\ : InMux
    port map (
            O => \N__55510\,
            I => \N__55507\
        );

    \I__13169\ : LocalMux
    port map (
            O => \N__55507\,
            I => \N__55504\
        );

    \I__13168\ : Odrv12
    port map (
            O => \N__55504\,
            I => n23348
        );

    \I__13167\ : InMux
    port map (
            O => \N__55501\,
            I => \N__55498\
        );

    \I__13166\ : LocalMux
    port map (
            O => \N__55498\,
            I => \N__55494\
        );

    \I__13165\ : CascadeMux
    port map (
            O => \N__55497\,
            I => \N__55491\
        );

    \I__13164\ : Span4Mux_h
    port map (
            O => \N__55494\,
            I => \N__55487\
        );

    \I__13163\ : InMux
    port map (
            O => \N__55491\,
            I => \N__55482\
        );

    \I__13162\ : InMux
    port map (
            O => \N__55490\,
            I => \N__55482\
        );

    \I__13161\ : Odrv4
    port map (
            O => \N__55487\,
            I => req_data_cnt_7
        );

    \I__13160\ : LocalMux
    port map (
            O => \N__55482\,
            I => req_data_cnt_7
        );

    \I__13159\ : InMux
    port map (
            O => \N__55477\,
            I => \N__55474\
        );

    \I__13158\ : LocalMux
    port map (
            O => \N__55474\,
            I => \N__55471\
        );

    \I__13157\ : Span12Mux_v
    port map (
            O => \N__55471\,
            I => \N__55466\
        );

    \I__13156\ : InMux
    port map (
            O => \N__55470\,
            I => \N__55461\
        );

    \I__13155\ : InMux
    port map (
            O => \N__55469\,
            I => \N__55461\
        );

    \I__13154\ : Odrv12
    port map (
            O => \N__55466\,
            I => \acadc_skipCount_7\
        );

    \I__13153\ : LocalMux
    port map (
            O => \N__55461\,
            I => \acadc_skipCount_7\
        );

    \I__13152\ : InMux
    port map (
            O => \N__55456\,
            I => \N__55453\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__55453\,
            I => n22262
        );

    \I__13150\ : InMux
    port map (
            O => \N__55450\,
            I => \N__55447\
        );

    \I__13149\ : LocalMux
    port map (
            O => \N__55447\,
            I => \N__55444\
        );

    \I__13148\ : Odrv12
    port map (
            O => \N__55444\,
            I => buf_data_iac_14
        );

    \I__13147\ : InMux
    port map (
            O => \N__55441\,
            I => \N__55438\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__55438\,
            I => \N__55435\
        );

    \I__13145\ : Odrv4
    port map (
            O => \N__55435\,
            I => n22391
        );

    \I__13144\ : InMux
    port map (
            O => \N__55432\,
            I => \N__55427\
        );

    \I__13143\ : InMux
    port map (
            O => \N__55431\,
            I => \N__55424\
        );

    \I__13142\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55420\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__55427\,
            I => \N__55415\
        );

    \I__13140\ : LocalMux
    port map (
            O => \N__55424\,
            I => \N__55415\
        );

    \I__13139\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55412\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__55420\,
            I => \N__55409\
        );

    \I__13137\ : Span4Mux_v
    port map (
            O => \N__55415\,
            I => \N__55404\
        );

    \I__13136\ : LocalMux
    port map (
            O => \N__55412\,
            I => \N__55404\
        );

    \I__13135\ : Span4Mux_v
    port map (
            O => \N__55409\,
            I => \N__55394\
        );

    \I__13134\ : Span4Mux_v
    port map (
            O => \N__55404\,
            I => \N__55394\
        );

    \I__13133\ : InMux
    port map (
            O => \N__55403\,
            I => \N__55389\
        );

    \I__13132\ : InMux
    port map (
            O => \N__55402\,
            I => \N__55389\
        );

    \I__13131\ : InMux
    port map (
            O => \N__55401\,
            I => \N__55385\
        );

    \I__13130\ : CascadeMux
    port map (
            O => \N__55400\,
            I => \N__55382\
        );

    \I__13129\ : InMux
    port map (
            O => \N__55399\,
            I => \N__55377\
        );

    \I__13128\ : Span4Mux_h
    port map (
            O => \N__55394\,
            I => \N__55372\
        );

    \I__13127\ : LocalMux
    port map (
            O => \N__55389\,
            I => \N__55372\
        );

    \I__13126\ : InMux
    port map (
            O => \N__55388\,
            I => \N__55365\
        );

    \I__13125\ : LocalMux
    port map (
            O => \N__55385\,
            I => \N__55362\
        );

    \I__13124\ : InMux
    port map (
            O => \N__55382\,
            I => \N__55359\
        );

    \I__13123\ : InMux
    port map (
            O => \N__55381\,
            I => \N__55356\
        );

    \I__13122\ : InMux
    port map (
            O => \N__55380\,
            I => \N__55353\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__55377\,
            I => \N__55348\
        );

    \I__13120\ : Span4Mux_v
    port map (
            O => \N__55372\,
            I => \N__55348\
        );

    \I__13119\ : InMux
    port map (
            O => \N__55371\,
            I => \N__55345\
        );

    \I__13118\ : InMux
    port map (
            O => \N__55370\,
            I => \N__55338\
        );

    \I__13117\ : InMux
    port map (
            O => \N__55369\,
            I => \N__55338\
        );

    \I__13116\ : InMux
    port map (
            O => \N__55368\,
            I => \N__55338\
        );

    \I__13115\ : LocalMux
    port map (
            O => \N__55365\,
            I => \N__55335\
        );

    \I__13114\ : Span4Mux_h
    port map (
            O => \N__55362\,
            I => \N__55332\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__55359\,
            I => \N__55329\
        );

    \I__13112\ : LocalMux
    port map (
            O => \N__55356\,
            I => \N__55326\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__55353\,
            I => \N__55323\
        );

    \I__13110\ : Span4Mux_h
    port map (
            O => \N__55348\,
            I => \N__55320\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__55345\,
            I => \N__55313\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__55338\,
            I => \N__55313\
        );

    \I__13107\ : Sp12to4
    port map (
            O => \N__55335\,
            I => \N__55313\
        );

    \I__13106\ : Span4Mux_h
    port map (
            O => \N__55332\,
            I => \N__55310\
        );

    \I__13105\ : Span12Mux_h
    port map (
            O => \N__55329\,
            I => \N__55307\
        );

    \I__13104\ : Span4Mux_v
    port map (
            O => \N__55326\,
            I => \N__55304\
        );

    \I__13103\ : Span12Mux_v
    port map (
            O => \N__55323\,
            I => \N__55297\
        );

    \I__13102\ : Sp12to4
    port map (
            O => \N__55320\,
            I => \N__55297\
        );

    \I__13101\ : Span12Mux_v
    port map (
            O => \N__55313\,
            I => \N__55297\
        );

    \I__13100\ : Odrv4
    port map (
            O => \N__55310\,
            I => n12509
        );

    \I__13099\ : Odrv12
    port map (
            O => \N__55307\,
            I => n12509
        );

    \I__13098\ : Odrv4
    port map (
            O => \N__55304\,
            I => n12509
        );

    \I__13097\ : Odrv12
    port map (
            O => \N__55297\,
            I => n12509
        );

    \I__13096\ : InMux
    port map (
            O => \N__55288\,
            I => \N__55284\
        );

    \I__13095\ : InMux
    port map (
            O => \N__55287\,
            I => \N__55280\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__55284\,
            I => \N__55277\
        );

    \I__13093\ : CascadeMux
    port map (
            O => \N__55283\,
            I => \N__55273\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__55280\,
            I => \N__55270\
        );

    \I__13091\ : Sp12to4
    port map (
            O => \N__55277\,
            I => \N__55267\
        );

    \I__13090\ : InMux
    port map (
            O => \N__55276\,
            I => \N__55264\
        );

    \I__13089\ : InMux
    port map (
            O => \N__55273\,
            I => \N__55261\
        );

    \I__13088\ : Span4Mux_v
    port map (
            O => \N__55270\,
            I => \N__55258\
        );

    \I__13087\ : Span12Mux_v
    port map (
            O => \N__55267\,
            I => \N__55255\
        );

    \I__13086\ : LocalMux
    port map (
            O => \N__55264\,
            I => \N__55252\
        );

    \I__13085\ : LocalMux
    port map (
            O => \N__55261\,
            I => \N__55249\
        );

    \I__13084\ : Span4Mux_h
    port map (
            O => \N__55258\,
            I => \N__55246\
        );

    \I__13083\ : Odrv12
    port map (
            O => \N__55255\,
            I => n14_adj_1660
        );

    \I__13082\ : Odrv4
    port map (
            O => \N__55252\,
            I => n14_adj_1660
        );

    \I__13081\ : Odrv4
    port map (
            O => \N__55249\,
            I => n14_adj_1660
        );

    \I__13080\ : Odrv4
    port map (
            O => \N__55246\,
            I => n14_adj_1660
        );

    \I__13079\ : InMux
    port map (
            O => \N__55237\,
            I => \N__55234\
        );

    \I__13078\ : LocalMux
    port map (
            O => \N__55234\,
            I => \N__55231\
        );

    \I__13077\ : Span4Mux_v
    port map (
            O => \N__55231\,
            I => \N__55228\
        );

    \I__13076\ : Sp12to4
    port map (
            O => \N__55228\,
            I => \N__55224\
        );

    \I__13075\ : InMux
    port map (
            O => \N__55227\,
            I => \N__55220\
        );

    \I__13074\ : Span12Mux_h
    port map (
            O => \N__55224\,
            I => \N__55217\
        );

    \I__13073\ : InMux
    port map (
            O => \N__55223\,
            I => \N__55214\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__55220\,
            I => buf_dds1_13
        );

    \I__13071\ : Odrv12
    port map (
            O => \N__55217\,
            I => buf_dds1_13
        );

    \I__13070\ : LocalMux
    port map (
            O => \N__55214\,
            I => buf_dds1_13
        );

    \I__13069\ : InMux
    port map (
            O => \N__55207\,
            I => \N__55203\
        );

    \I__13068\ : InMux
    port map (
            O => \N__55206\,
            I => \N__55200\
        );

    \I__13067\ : LocalMux
    port map (
            O => \N__55203\,
            I => \N__55195\
        );

    \I__13066\ : LocalMux
    port map (
            O => \N__55200\,
            I => \N__55195\
        );

    \I__13065\ : Span4Mux_v
    port map (
            O => \N__55195\,
            I => \N__55190\
        );

    \I__13064\ : CascadeMux
    port map (
            O => \N__55194\,
            I => \N__55186\
        );

    \I__13063\ : CascadeMux
    port map (
            O => \N__55193\,
            I => \N__55183\
        );

    \I__13062\ : Span4Mux_h
    port map (
            O => \N__55190\,
            I => \N__55180\
        );

    \I__13061\ : InMux
    port map (
            O => \N__55189\,
            I => \N__55177\
        );

    \I__13060\ : InMux
    port map (
            O => \N__55186\,
            I => \N__55174\
        );

    \I__13059\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55171\
        );

    \I__13058\ : Span4Mux_v
    port map (
            O => \N__55180\,
            I => \N__55164\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__55177\,
            I => \N__55164\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__55174\,
            I => \N__55161\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__55171\,
            I => \N__55157\
        );

    \I__13054\ : InMux
    port map (
            O => \N__55170\,
            I => \N__55154\
        );

    \I__13053\ : CascadeMux
    port map (
            O => \N__55169\,
            I => \N__55151\
        );

    \I__13052\ : Span4Mux_v
    port map (
            O => \N__55164\,
            I => \N__55148\
        );

    \I__13051\ : Span4Mux_v
    port map (
            O => \N__55161\,
            I => \N__55145\
        );

    \I__13050\ : InMux
    port map (
            O => \N__55160\,
            I => \N__55142\
        );

    \I__13049\ : Span4Mux_v
    port map (
            O => \N__55157\,
            I => \N__55139\
        );

    \I__13048\ : LocalMux
    port map (
            O => \N__55154\,
            I => \N__55136\
        );

    \I__13047\ : InMux
    port map (
            O => \N__55151\,
            I => \N__55133\
        );

    \I__13046\ : Span4Mux_h
    port map (
            O => \N__55148\,
            I => \N__55129\
        );

    \I__13045\ : Sp12to4
    port map (
            O => \N__55145\,
            I => \N__55124\
        );

    \I__13044\ : LocalMux
    port map (
            O => \N__55142\,
            I => \N__55124\
        );

    \I__13043\ : Span4Mux_h
    port map (
            O => \N__55139\,
            I => \N__55117\
        );

    \I__13042\ : Span4Mux_h
    port map (
            O => \N__55136\,
            I => \N__55117\
        );

    \I__13041\ : LocalMux
    port map (
            O => \N__55133\,
            I => \N__55117\
        );

    \I__13040\ : InMux
    port map (
            O => \N__55132\,
            I => \N__55114\
        );

    \I__13039\ : Odrv4
    port map (
            O => \N__55129\,
            I => comm_rx_buf_5
        );

    \I__13038\ : Odrv12
    port map (
            O => \N__55124\,
            I => comm_rx_buf_5
        );

    \I__13037\ : Odrv4
    port map (
            O => \N__55117\,
            I => comm_rx_buf_5
        );

    \I__13036\ : LocalMux
    port map (
            O => \N__55114\,
            I => comm_rx_buf_5
        );

    \I__13035\ : InMux
    port map (
            O => \N__55105\,
            I => \N__55102\
        );

    \I__13034\ : LocalMux
    port map (
            O => \N__55102\,
            I => \N__55099\
        );

    \I__13033\ : Span4Mux_h
    port map (
            O => \N__55099\,
            I => \N__55096\
        );

    \I__13032\ : Odrv4
    port map (
            O => \N__55096\,
            I => buf_data_vac_13
        );

    \I__13031\ : InMux
    port map (
            O => \N__55093\,
            I => \N__55090\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__55090\,
            I => \N__55087\
        );

    \I__13029\ : Span4Mux_h
    port map (
            O => \N__55087\,
            I => \N__55084\
        );

    \I__13028\ : Odrv4
    port map (
            O => \N__55084\,
            I => comm_buf_4_5
        );

    \I__13027\ : CascadeMux
    port map (
            O => \N__55081\,
            I => \N__55078\
        );

    \I__13026\ : InMux
    port map (
            O => \N__55078\,
            I => \N__55073\
        );

    \I__13025\ : InMux
    port map (
            O => \N__55077\,
            I => \N__55068\
        );

    \I__13024\ : CascadeMux
    port map (
            O => \N__55076\,
            I => \N__55064\
        );

    \I__13023\ : LocalMux
    port map (
            O => \N__55073\,
            I => \N__55061\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55072\,
            I => \N__55057\
        );

    \I__13021\ : InMux
    port map (
            O => \N__55071\,
            I => \N__55054\
        );

    \I__13020\ : LocalMux
    port map (
            O => \N__55068\,
            I => \N__55051\
        );

    \I__13019\ : InMux
    port map (
            O => \N__55067\,
            I => \N__55048\
        );

    \I__13018\ : InMux
    port map (
            O => \N__55064\,
            I => \N__55045\
        );

    \I__13017\ : Span4Mux_v
    port map (
            O => \N__55061\,
            I => \N__55042\
        );

    \I__13016\ : InMux
    port map (
            O => \N__55060\,
            I => \N__55039\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__55057\,
            I => \N__55033\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__55054\,
            I => \N__55033\
        );

    \I__13013\ : Span4Mux_v
    port map (
            O => \N__55051\,
            I => \N__55028\
        );

    \I__13012\ : LocalMux
    port map (
            O => \N__55048\,
            I => \N__55028\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__55045\,
            I => \N__55025\
        );

    \I__13010\ : Span4Mux_h
    port map (
            O => \N__55042\,
            I => \N__55020\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__55039\,
            I => \N__55020\
        );

    \I__13008\ : InMux
    port map (
            O => \N__55038\,
            I => \N__55017\
        );

    \I__13007\ : Span12Mux_v
    port map (
            O => \N__55033\,
            I => \N__55013\
        );

    \I__13006\ : Span4Mux_h
    port map (
            O => \N__55028\,
            I => \N__55010\
        );

    \I__13005\ : Span12Mux_h
    port map (
            O => \N__55025\,
            I => \N__55003\
        );

    \I__13004\ : Sp12to4
    port map (
            O => \N__55020\,
            I => \N__55003\
        );

    \I__13003\ : LocalMux
    port map (
            O => \N__55017\,
            I => \N__55003\
        );

    \I__13002\ : InMux
    port map (
            O => \N__55016\,
            I => \N__55000\
        );

    \I__13001\ : Odrv12
    port map (
            O => \N__55013\,
            I => comm_rx_buf_4
        );

    \I__13000\ : Odrv4
    port map (
            O => \N__55010\,
            I => comm_rx_buf_4
        );

    \I__12999\ : Odrv12
    port map (
            O => \N__55003\,
            I => comm_rx_buf_4
        );

    \I__12998\ : LocalMux
    port map (
            O => \N__55000\,
            I => comm_rx_buf_4
        );

    \I__12997\ : InMux
    port map (
            O => \N__54991\,
            I => \N__54988\
        );

    \I__12996\ : LocalMux
    port map (
            O => \N__54988\,
            I => \N__54985\
        );

    \I__12995\ : Span12Mux_v
    port map (
            O => \N__54985\,
            I => \N__54982\
        );

    \I__12994\ : Odrv12
    port map (
            O => \N__54982\,
            I => buf_data_vac_12
        );

    \I__12993\ : InMux
    port map (
            O => \N__54979\,
            I => \N__54976\
        );

    \I__12992\ : LocalMux
    port map (
            O => \N__54976\,
            I => \N__54973\
        );

    \I__12991\ : Span4Mux_v
    port map (
            O => \N__54973\,
            I => \N__54970\
        );

    \I__12990\ : Span4Mux_h
    port map (
            O => \N__54970\,
            I => \N__54967\
        );

    \I__12989\ : Odrv4
    port map (
            O => \N__54967\,
            I => comm_buf_4_4
        );

    \I__12988\ : InMux
    port map (
            O => \N__54964\,
            I => \N__54961\
        );

    \I__12987\ : LocalMux
    port map (
            O => \N__54961\,
            I => \N__54958\
        );

    \I__12986\ : Span4Mux_h
    port map (
            O => \N__54958\,
            I => \N__54955\
        );

    \I__12985\ : Span4Mux_v
    port map (
            O => \N__54955\,
            I => \N__54952\
        );

    \I__12984\ : Odrv4
    port map (
            O => \N__54952\,
            I => buf_data_vac_11
        );

    \I__12983\ : InMux
    port map (
            O => \N__54949\,
            I => \N__54946\
        );

    \I__12982\ : LocalMux
    port map (
            O => \N__54946\,
            I => \N__54943\
        );

    \I__12981\ : Odrv4
    port map (
            O => \N__54943\,
            I => comm_buf_4_3
        );

    \I__12980\ : InMux
    port map (
            O => \N__54940\,
            I => \N__54935\
        );

    \I__12979\ : InMux
    port map (
            O => \N__54939\,
            I => \N__54932\
        );

    \I__12978\ : InMux
    port map (
            O => \N__54938\,
            I => \N__54926\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__54935\,
            I => \N__54920\
        );

    \I__12976\ : LocalMux
    port map (
            O => \N__54932\,
            I => \N__54920\
        );

    \I__12975\ : InMux
    port map (
            O => \N__54931\,
            I => \N__54917\
        );

    \I__12974\ : InMux
    port map (
            O => \N__54930\,
            I => \N__54914\
        );

    \I__12973\ : InMux
    port map (
            O => \N__54929\,
            I => \N__54911\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__54926\,
            I => \N__54908\
        );

    \I__12971\ : InMux
    port map (
            O => \N__54925\,
            I => \N__54905\
        );

    \I__12970\ : Span4Mux_v
    port map (
            O => \N__54920\,
            I => \N__54900\
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__54917\,
            I => \N__54900\
        );

    \I__12968\ : LocalMux
    port map (
            O => \N__54914\,
            I => \N__54897\
        );

    \I__12967\ : LocalMux
    port map (
            O => \N__54911\,
            I => \N__54893\
        );

    \I__12966\ : Span4Mux_v
    port map (
            O => \N__54908\,
            I => \N__54888\
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__54905\,
            I => \N__54888\
        );

    \I__12964\ : Span4Mux_h
    port map (
            O => \N__54900\,
            I => \N__54885\
        );

    \I__12963\ : Span4Mux_v
    port map (
            O => \N__54897\,
            I => \N__54882\
        );

    \I__12962\ : InMux
    port map (
            O => \N__54896\,
            I => \N__54879\
        );

    \I__12961\ : Span12Mux_v
    port map (
            O => \N__54893\,
            I => \N__54875\
        );

    \I__12960\ : Span4Mux_h
    port map (
            O => \N__54888\,
            I => \N__54872\
        );

    \I__12959\ : Span4Mux_v
    port map (
            O => \N__54885\,
            I => \N__54869\
        );

    \I__12958\ : Span4Mux_h
    port map (
            O => \N__54882\,
            I => \N__54864\
        );

    \I__12957\ : LocalMux
    port map (
            O => \N__54879\,
            I => \N__54864\
        );

    \I__12956\ : InMux
    port map (
            O => \N__54878\,
            I => \N__54861\
        );

    \I__12955\ : Odrv12
    port map (
            O => \N__54875\,
            I => comm_rx_buf_2
        );

    \I__12954\ : Odrv4
    port map (
            O => \N__54872\,
            I => comm_rx_buf_2
        );

    \I__12953\ : Odrv4
    port map (
            O => \N__54869\,
            I => comm_rx_buf_2
        );

    \I__12952\ : Odrv4
    port map (
            O => \N__54864\,
            I => comm_rx_buf_2
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__54861\,
            I => comm_rx_buf_2
        );

    \I__12950\ : InMux
    port map (
            O => \N__54850\,
            I => \N__54847\
        );

    \I__12949\ : LocalMux
    port map (
            O => \N__54847\,
            I => \N__54844\
        );

    \I__12948\ : Span12Mux_v
    port map (
            O => \N__54844\,
            I => \N__54841\
        );

    \I__12947\ : Odrv12
    port map (
            O => \N__54841\,
            I => buf_data_vac_10
        );

    \I__12946\ : InMux
    port map (
            O => \N__54838\,
            I => \N__54835\
        );

    \I__12945\ : LocalMux
    port map (
            O => \N__54835\,
            I => \N__54832\
        );

    \I__12944\ : Span4Mux_h
    port map (
            O => \N__54832\,
            I => \N__54829\
        );

    \I__12943\ : Span4Mux_h
    port map (
            O => \N__54829\,
            I => \N__54826\
        );

    \I__12942\ : Odrv4
    port map (
            O => \N__54826\,
            I => comm_buf_4_2
        );

    \I__12941\ : CascadeMux
    port map (
            O => \N__54823\,
            I => \N__54820\
        );

    \I__12940\ : InMux
    port map (
            O => \N__54820\,
            I => \N__54817\
        );

    \I__12939\ : LocalMux
    port map (
            O => \N__54817\,
            I => \N__54813\
        );

    \I__12938\ : InMux
    port map (
            O => \N__54816\,
            I => \N__54810\
        );

    \I__12937\ : Span4Mux_v
    port map (
            O => \N__54813\,
            I => \N__54804\
        );

    \I__12936\ : LocalMux
    port map (
            O => \N__54810\,
            I => \N__54804\
        );

    \I__12935\ : InMux
    port map (
            O => \N__54809\,
            I => \N__54801\
        );

    \I__12934\ : Span4Mux_v
    port map (
            O => \N__54804\,
            I => \N__54797\
        );

    \I__12933\ : LocalMux
    port map (
            O => \N__54801\,
            I => \N__54793\
        );

    \I__12932\ : InMux
    port map (
            O => \N__54800\,
            I => \N__54789\
        );

    \I__12931\ : Span4Mux_h
    port map (
            O => \N__54797\,
            I => \N__54785\
        );

    \I__12930\ : InMux
    port map (
            O => \N__54796\,
            I => \N__54782\
        );

    \I__12929\ : Span4Mux_h
    port map (
            O => \N__54793\,
            I => \N__54779\
        );

    \I__12928\ : InMux
    port map (
            O => \N__54792\,
            I => \N__54776\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__54789\,
            I => \N__54773\
        );

    \I__12926\ : InMux
    port map (
            O => \N__54788\,
            I => \N__54770\
        );

    \I__12925\ : Span4Mux_h
    port map (
            O => \N__54785\,
            I => \N__54764\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__54782\,
            I => \N__54764\
        );

    \I__12923\ : Span4Mux_v
    port map (
            O => \N__54779\,
            I => \N__54759\
        );

    \I__12922\ : LocalMux
    port map (
            O => \N__54776\,
            I => \N__54759\
        );

    \I__12921\ : Span4Mux_v
    port map (
            O => \N__54773\,
            I => \N__54754\
        );

    \I__12920\ : LocalMux
    port map (
            O => \N__54770\,
            I => \N__54754\
        );

    \I__12919\ : InMux
    port map (
            O => \N__54769\,
            I => \N__54751\
        );

    \I__12918\ : Span4Mux_v
    port map (
            O => \N__54764\,
            I => \N__54747\
        );

    \I__12917\ : Span4Mux_h
    port map (
            O => \N__54759\,
            I => \N__54744\
        );

    \I__12916\ : Span4Mux_h
    port map (
            O => \N__54754\,
            I => \N__54741\
        );

    \I__12915\ : LocalMux
    port map (
            O => \N__54751\,
            I => \N__54738\
        );

    \I__12914\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54735\
        );

    \I__12913\ : Odrv4
    port map (
            O => \N__54747\,
            I => comm_rx_buf_1
        );

    \I__12912\ : Odrv4
    port map (
            O => \N__54744\,
            I => comm_rx_buf_1
        );

    \I__12911\ : Odrv4
    port map (
            O => \N__54741\,
            I => comm_rx_buf_1
        );

    \I__12910\ : Odrv4
    port map (
            O => \N__54738\,
            I => comm_rx_buf_1
        );

    \I__12909\ : LocalMux
    port map (
            O => \N__54735\,
            I => comm_rx_buf_1
        );

    \I__12908\ : InMux
    port map (
            O => \N__54724\,
            I => \N__54721\
        );

    \I__12907\ : LocalMux
    port map (
            O => \N__54721\,
            I => \N__54718\
        );

    \I__12906\ : Span4Mux_h
    port map (
            O => \N__54718\,
            I => \N__54715\
        );

    \I__12905\ : Span4Mux_v
    port map (
            O => \N__54715\,
            I => \N__54712\
        );

    \I__12904\ : Odrv4
    port map (
            O => \N__54712\,
            I => buf_data_vac_9
        );

    \I__12903\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54706\
        );

    \I__12902\ : LocalMux
    port map (
            O => \N__54706\,
            I => \N__54703\
        );

    \I__12901\ : Span4Mux_h
    port map (
            O => \N__54703\,
            I => \N__54700\
        );

    \I__12900\ : Span4Mux_v
    port map (
            O => \N__54700\,
            I => \N__54697\
        );

    \I__12899\ : Odrv4
    port map (
            O => \N__54697\,
            I => comm_buf_4_1
        );

    \I__12898\ : CEMux
    port map (
            O => \N__54694\,
            I => \N__54691\
        );

    \I__12897\ : LocalMux
    port map (
            O => \N__54691\,
            I => n12892
        );

    \I__12896\ : SRMux
    port map (
            O => \N__54688\,
            I => \N__54685\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__54685\,
            I => \N__54682\
        );

    \I__12894\ : Span4Mux_h
    port map (
            O => \N__54682\,
            I => \N__54679\
        );

    \I__12893\ : Odrv4
    port map (
            O => \N__54679\,
            I => n15510
        );

    \I__12892\ : InMux
    port map (
            O => \N__54676\,
            I => \N__54673\
        );

    \I__12891\ : LocalMux
    port map (
            O => \N__54673\,
            I => \N__54669\
        );

    \I__12890\ : InMux
    port map (
            O => \N__54672\,
            I => \N__54666\
        );

    \I__12889\ : Span4Mux_h
    port map (
            O => \N__54669\,
            I => \N__54663\
        );

    \I__12888\ : LocalMux
    port map (
            O => \N__54666\,
            I => data_idxvec_7
        );

    \I__12887\ : Odrv4
    port map (
            O => \N__54663\,
            I => data_idxvec_7
        );

    \I__12886\ : InMux
    port map (
            O => \N__54658\,
            I => \N__54654\
        );

    \I__12885\ : InMux
    port map (
            O => \N__54657\,
            I => \N__54651\
        );

    \I__12884\ : LocalMux
    port map (
            O => \N__54654\,
            I => \N__54647\
        );

    \I__12883\ : LocalMux
    port map (
            O => \N__54651\,
            I => \N__54644\
        );

    \I__12882\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54641\
        );

    \I__12881\ : Span4Mux_h
    port map (
            O => \N__54647\,
            I => \N__54638\
        );

    \I__12880\ : Span4Mux_h
    port map (
            O => \N__54644\,
            I => \N__54635\
        );

    \I__12879\ : LocalMux
    port map (
            O => \N__54641\,
            I => data_cntvec_7
        );

    \I__12878\ : Odrv4
    port map (
            O => \N__54638\,
            I => data_cntvec_7
        );

    \I__12877\ : Odrv4
    port map (
            O => \N__54635\,
            I => data_cntvec_7
        );

    \I__12876\ : InMux
    port map (
            O => \N__54628\,
            I => \N__54625\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__54625\,
            I => \N__54622\
        );

    \I__12874\ : Odrv12
    port map (
            O => \N__54622\,
            I => buf_data_iac_15
        );

    \I__12873\ : CascadeMux
    port map (
            O => \N__54619\,
            I => \n26_adj_1716_cascade_\
        );

    \I__12872\ : CascadeMux
    port map (
            O => \N__54616\,
            I => \n22263_cascade_\
        );

    \I__12871\ : InMux
    port map (
            O => \N__54613\,
            I => \N__54603\
        );

    \I__12870\ : InMux
    port map (
            O => \N__54612\,
            I => \N__54603\
        );

    \I__12869\ : InMux
    port map (
            O => \N__54611\,
            I => \N__54596\
        );

    \I__12868\ : InMux
    port map (
            O => \N__54610\,
            I => \N__54593\
        );

    \I__12867\ : InMux
    port map (
            O => \N__54609\,
            I => \N__54590\
        );

    \I__12866\ : InMux
    port map (
            O => \N__54608\,
            I => \N__54581\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__54603\,
            I => \N__54578\
        );

    \I__12864\ : InMux
    port map (
            O => \N__54602\,
            I => \N__54573\
        );

    \I__12863\ : InMux
    port map (
            O => \N__54601\,
            I => \N__54573\
        );

    \I__12862\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54567\
        );

    \I__12861\ : InMux
    port map (
            O => \N__54599\,
            I => \N__54567\
        );

    \I__12860\ : LocalMux
    port map (
            O => \N__54596\,
            I => \N__54562\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__54593\,
            I => \N__54562\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__54590\,
            I => \N__54559\
        );

    \I__12857\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54550\
        );

    \I__12856\ : InMux
    port map (
            O => \N__54588\,
            I => \N__54550\
        );

    \I__12855\ : InMux
    port map (
            O => \N__54587\,
            I => \N__54550\
        );

    \I__12854\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54550\
        );

    \I__12853\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54547\
        );

    \I__12852\ : InMux
    port map (
            O => \N__54584\,
            I => \N__54543\
        );

    \I__12851\ : LocalMux
    port map (
            O => \N__54581\,
            I => \N__54534\
        );

    \I__12850\ : Span4Mux_h
    port map (
            O => \N__54578\,
            I => \N__54529\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__54573\,
            I => \N__54529\
        );

    \I__12848\ : InMux
    port map (
            O => \N__54572\,
            I => \N__54522\
        );

    \I__12847\ : LocalMux
    port map (
            O => \N__54567\,
            I => \N__54513\
        );

    \I__12846\ : Span4Mux_v
    port map (
            O => \N__54562\,
            I => \N__54513\
        );

    \I__12845\ : Span4Mux_v
    port map (
            O => \N__54559\,
            I => \N__54513\
        );

    \I__12844\ : LocalMux
    port map (
            O => \N__54550\,
            I => \N__54513\
        );

    \I__12843\ : LocalMux
    port map (
            O => \N__54547\,
            I => \N__54510\
        );

    \I__12842\ : InMux
    port map (
            O => \N__54546\,
            I => \N__54507\
        );

    \I__12841\ : LocalMux
    port map (
            O => \N__54543\,
            I => \N__54504\
        );

    \I__12840\ : InMux
    port map (
            O => \N__54542\,
            I => \N__54495\
        );

    \I__12839\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54495\
        );

    \I__12838\ : InMux
    port map (
            O => \N__54540\,
            I => \N__54495\
        );

    \I__12837\ : InMux
    port map (
            O => \N__54539\,
            I => \N__54495\
        );

    \I__12836\ : InMux
    port map (
            O => \N__54538\,
            I => \N__54490\
        );

    \I__12835\ : InMux
    port map (
            O => \N__54537\,
            I => \N__54490\
        );

    \I__12834\ : Span4Mux_h
    port map (
            O => \N__54534\,
            I => \N__54487\
        );

    \I__12833\ : Span4Mux_h
    port map (
            O => \N__54529\,
            I => \N__54484\
        );

    \I__12832\ : InMux
    port map (
            O => \N__54528\,
            I => \N__54475\
        );

    \I__12831\ : InMux
    port map (
            O => \N__54527\,
            I => \N__54475\
        );

    \I__12830\ : InMux
    port map (
            O => \N__54526\,
            I => \N__54475\
        );

    \I__12829\ : InMux
    port map (
            O => \N__54525\,
            I => \N__54475\
        );

    \I__12828\ : LocalMux
    port map (
            O => \N__54522\,
            I => \N__54468\
        );

    \I__12827\ : Span4Mux_h
    port map (
            O => \N__54513\,
            I => \N__54468\
        );

    \I__12826\ : Span4Mux_v
    port map (
            O => \N__54510\,
            I => \N__54468\
        );

    \I__12825\ : LocalMux
    port map (
            O => \N__54507\,
            I => \N__54465\
        );

    \I__12824\ : Span4Mux_h
    port map (
            O => \N__54504\,
            I => \N__54458\
        );

    \I__12823\ : LocalMux
    port map (
            O => \N__54495\,
            I => \N__54458\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__54490\,
            I => \N__54458\
        );

    \I__12821\ : Odrv4
    port map (
            O => \N__54487\,
            I => comm_index_2
        );

    \I__12820\ : Odrv4
    port map (
            O => \N__54484\,
            I => comm_index_2
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__54475\,
            I => comm_index_2
        );

    \I__12818\ : Odrv4
    port map (
            O => \N__54468\,
            I => comm_index_2
        );

    \I__12817\ : Odrv4
    port map (
            O => \N__54465\,
            I => comm_index_2
        );

    \I__12816\ : Odrv4
    port map (
            O => \N__54458\,
            I => comm_index_2
        );

    \I__12815\ : CascadeMux
    port map (
            O => \N__54445\,
            I => \N__54441\
        );

    \I__12814\ : InMux
    port map (
            O => \N__54444\,
            I => \N__54438\
        );

    \I__12813\ : InMux
    port map (
            O => \N__54441\,
            I => \N__54435\
        );

    \I__12812\ : LocalMux
    port map (
            O => \N__54438\,
            I => n21956
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__54435\,
            I => n21956
        );

    \I__12810\ : InMux
    port map (
            O => \N__54430\,
            I => \N__54427\
        );

    \I__12809\ : LocalMux
    port map (
            O => \N__54427\,
            I => n21862
        );

    \I__12808\ : CascadeMux
    port map (
            O => \N__54424\,
            I => \N__54410\
        );

    \I__12807\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54402\
        );

    \I__12806\ : InMux
    port map (
            O => \N__54422\,
            I => \N__54391\
        );

    \I__12805\ : InMux
    port map (
            O => \N__54421\,
            I => \N__54391\
        );

    \I__12804\ : InMux
    port map (
            O => \N__54420\,
            I => \N__54391\
        );

    \I__12803\ : InMux
    port map (
            O => \N__54419\,
            I => \N__54388\
        );

    \I__12802\ : CascadeMux
    port map (
            O => \N__54418\,
            I => \N__54385\
        );

    \I__12801\ : CascadeMux
    port map (
            O => \N__54417\,
            I => \N__54382\
        );

    \I__12800\ : InMux
    port map (
            O => \N__54416\,
            I => \N__54373\
        );

    \I__12799\ : InMux
    port map (
            O => \N__54415\,
            I => \N__54373\
        );

    \I__12798\ : InMux
    port map (
            O => \N__54414\,
            I => \N__54373\
        );

    \I__12797\ : InMux
    port map (
            O => \N__54413\,
            I => \N__54373\
        );

    \I__12796\ : InMux
    port map (
            O => \N__54410\,
            I => \N__54367\
        );

    \I__12795\ : InMux
    port map (
            O => \N__54409\,
            I => \N__54364\
        );

    \I__12794\ : InMux
    port map (
            O => \N__54408\,
            I => \N__54353\
        );

    \I__12793\ : InMux
    port map (
            O => \N__54407\,
            I => \N__54353\
        );

    \I__12792\ : InMux
    port map (
            O => \N__54406\,
            I => \N__54353\
        );

    \I__12791\ : InMux
    port map (
            O => \N__54405\,
            I => \N__54353\
        );

    \I__12790\ : LocalMux
    port map (
            O => \N__54402\,
            I => \N__54350\
        );

    \I__12789\ : InMux
    port map (
            O => \N__54401\,
            I => \N__54341\
        );

    \I__12788\ : InMux
    port map (
            O => \N__54400\,
            I => \N__54341\
        );

    \I__12787\ : InMux
    port map (
            O => \N__54399\,
            I => \N__54341\
        );

    \I__12786\ : InMux
    port map (
            O => \N__54398\,
            I => \N__54341\
        );

    \I__12785\ : LocalMux
    port map (
            O => \N__54391\,
            I => \N__54338\
        );

    \I__12784\ : LocalMux
    port map (
            O => \N__54388\,
            I => \N__54335\
        );

    \I__12783\ : InMux
    port map (
            O => \N__54385\,
            I => \N__54332\
        );

    \I__12782\ : InMux
    port map (
            O => \N__54382\,
            I => \N__54327\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__54373\,
            I => \N__54323\
        );

    \I__12780\ : InMux
    port map (
            O => \N__54372\,
            I => \N__54316\
        );

    \I__12779\ : InMux
    port map (
            O => \N__54371\,
            I => \N__54316\
        );

    \I__12778\ : InMux
    port map (
            O => \N__54370\,
            I => \N__54316\
        );

    \I__12777\ : LocalMux
    port map (
            O => \N__54367\,
            I => \N__54313\
        );

    \I__12776\ : LocalMux
    port map (
            O => \N__54364\,
            I => \N__54303\
        );

    \I__12775\ : InMux
    port map (
            O => \N__54363\,
            I => \N__54298\
        );

    \I__12774\ : InMux
    port map (
            O => \N__54362\,
            I => \N__54298\
        );

    \I__12773\ : LocalMux
    port map (
            O => \N__54353\,
            I => \N__54293\
        );

    \I__12772\ : Span4Mux_v
    port map (
            O => \N__54350\,
            I => \N__54293\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__54341\,
            I => \N__54290\
        );

    \I__12770\ : Span4Mux_v
    port map (
            O => \N__54338\,
            I => \N__54287\
        );

    \I__12769\ : Span4Mux_h
    port map (
            O => \N__54335\,
            I => \N__54282\
        );

    \I__12768\ : LocalMux
    port map (
            O => \N__54332\,
            I => \N__54282\
        );

    \I__12767\ : InMux
    port map (
            O => \N__54331\,
            I => \N__54277\
        );

    \I__12766\ : InMux
    port map (
            O => \N__54330\,
            I => \N__54277\
        );

    \I__12765\ : LocalMux
    port map (
            O => \N__54327\,
            I => \N__54274\
        );

    \I__12764\ : InMux
    port map (
            O => \N__54326\,
            I => \N__54271\
        );

    \I__12763\ : Span4Mux_v
    port map (
            O => \N__54323\,
            I => \N__54264\
        );

    \I__12762\ : LocalMux
    port map (
            O => \N__54316\,
            I => \N__54264\
        );

    \I__12761\ : Span4Mux_h
    port map (
            O => \N__54313\,
            I => \N__54264\
        );

    \I__12760\ : InMux
    port map (
            O => \N__54312\,
            I => \N__54259\
        );

    \I__12759\ : InMux
    port map (
            O => \N__54311\,
            I => \N__54259\
        );

    \I__12758\ : InMux
    port map (
            O => \N__54310\,
            I => \N__54254\
        );

    \I__12757\ : InMux
    port map (
            O => \N__54309\,
            I => \N__54254\
        );

    \I__12756\ : InMux
    port map (
            O => \N__54308\,
            I => \N__54251\
        );

    \I__12755\ : InMux
    port map (
            O => \N__54307\,
            I => \N__54246\
        );

    \I__12754\ : InMux
    port map (
            O => \N__54306\,
            I => \N__54246\
        );

    \I__12753\ : Span4Mux_h
    port map (
            O => \N__54303\,
            I => \N__54243\
        );

    \I__12752\ : LocalMux
    port map (
            O => \N__54298\,
            I => \N__54234\
        );

    \I__12751\ : Span4Mux_h
    port map (
            O => \N__54293\,
            I => \N__54234\
        );

    \I__12750\ : Span4Mux_v
    port map (
            O => \N__54290\,
            I => \N__54234\
        );

    \I__12749\ : Span4Mux_h
    port map (
            O => \N__54287\,
            I => \N__54234\
        );

    \I__12748\ : Span4Mux_h
    port map (
            O => \N__54282\,
            I => \N__54231\
        );

    \I__12747\ : LocalMux
    port map (
            O => \N__54277\,
            I => \N__54220\
        );

    \I__12746\ : Span4Mux_h
    port map (
            O => \N__54274\,
            I => \N__54220\
        );

    \I__12745\ : LocalMux
    port map (
            O => \N__54271\,
            I => \N__54220\
        );

    \I__12744\ : Span4Mux_h
    port map (
            O => \N__54264\,
            I => \N__54220\
        );

    \I__12743\ : LocalMux
    port map (
            O => \N__54259\,
            I => \N__54220\
        );

    \I__12742\ : LocalMux
    port map (
            O => \N__54254\,
            I => comm_index_0
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__54251\,
            I => comm_index_0
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__54246\,
            I => comm_index_0
        );

    \I__12739\ : Odrv4
    port map (
            O => \N__54243\,
            I => comm_index_0
        );

    \I__12738\ : Odrv4
    port map (
            O => \N__54234\,
            I => comm_index_0
        );

    \I__12737\ : Odrv4
    port map (
            O => \N__54231\,
            I => comm_index_0
        );

    \I__12736\ : Odrv4
    port map (
            O => \N__54220\,
            I => comm_index_0
        );

    \I__12735\ : CascadeMux
    port map (
            O => \N__54205\,
            I => \n21862_cascade_\
        );

    \I__12734\ : InMux
    port map (
            O => \N__54202\,
            I => \N__54199\
        );

    \I__12733\ : LocalMux
    port map (
            O => \N__54199\,
            I => \N__54195\
        );

    \I__12732\ : InMux
    port map (
            O => \N__54198\,
            I => \N__54192\
        );

    \I__12731\ : Span4Mux_h
    port map (
            O => \N__54195\,
            I => \N__54189\
        );

    \I__12730\ : LocalMux
    port map (
            O => \N__54192\,
            I => n30_adj_1720
        );

    \I__12729\ : Odrv4
    port map (
            O => \N__54189\,
            I => n30_adj_1720
        );

    \I__12728\ : CascadeMux
    port map (
            O => \N__54184\,
            I => \N__54179\
        );

    \I__12727\ : CascadeMux
    port map (
            O => \N__54183\,
            I => \N__54176\
        );

    \I__12726\ : InMux
    port map (
            O => \N__54182\,
            I => \N__54172\
        );

    \I__12725\ : InMux
    port map (
            O => \N__54179\,
            I => \N__54168\
        );

    \I__12724\ : InMux
    port map (
            O => \N__54176\,
            I => \N__54165\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54175\,
            I => \N__54162\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__54172\,
            I => \N__54156\
        );

    \I__12721\ : InMux
    port map (
            O => \N__54171\,
            I => \N__54153\
        );

    \I__12720\ : LocalMux
    port map (
            O => \N__54168\,
            I => \N__54150\
        );

    \I__12719\ : LocalMux
    port map (
            O => \N__54165\,
            I => \N__54145\
        );

    \I__12718\ : LocalMux
    port map (
            O => \N__54162\,
            I => \N__54145\
        );

    \I__12717\ : CascadeMux
    port map (
            O => \N__54161\,
            I => \N__54142\
        );

    \I__12716\ : InMux
    port map (
            O => \N__54160\,
            I => \N__54137\
        );

    \I__12715\ : InMux
    port map (
            O => \N__54159\,
            I => \N__54137\
        );

    \I__12714\ : Span4Mux_h
    port map (
            O => \N__54156\,
            I => \N__54131\
        );

    \I__12713\ : LocalMux
    port map (
            O => \N__54153\,
            I => \N__54131\
        );

    \I__12712\ : Span4Mux_v
    port map (
            O => \N__54150\,
            I => \N__54128\
        );

    \I__12711\ : Span4Mux_h
    port map (
            O => \N__54145\,
            I => \N__54125\
        );

    \I__12710\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54122\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__54137\,
            I => \N__54119\
        );

    \I__12708\ : InMux
    port map (
            O => \N__54136\,
            I => \N__54116\
        );

    \I__12707\ : Span4Mux_h
    port map (
            O => \N__54131\,
            I => \N__54113\
        );

    \I__12706\ : Span4Mux_h
    port map (
            O => \N__54128\,
            I => \N__54110\
        );

    \I__12705\ : Span4Mux_v
    port map (
            O => \N__54125\,
            I => \N__54101\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__54122\,
            I => \N__54101\
        );

    \I__12703\ : Span4Mux_h
    port map (
            O => \N__54119\,
            I => \N__54101\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__54116\,
            I => \N__54101\
        );

    \I__12701\ : Span4Mux_v
    port map (
            O => \N__54113\,
            I => \N__54098\
        );

    \I__12700\ : Odrv4
    port map (
            O => \N__54110\,
            I => n21968
        );

    \I__12699\ : Odrv4
    port map (
            O => \N__54101\,
            I => n21968
        );

    \I__12698\ : Odrv4
    port map (
            O => \N__54098\,
            I => n21968
        );

    \I__12697\ : CascadeMux
    port map (
            O => \N__54091\,
            I => \n22_adj_1725_cascade_\
        );

    \I__12696\ : CascadeMux
    port map (
            O => \N__54088\,
            I => \n12677_cascade_\
        );

    \I__12695\ : InMux
    port map (
            O => \N__54085\,
            I => \N__54082\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__54082\,
            I => \N__54078\
        );

    \I__12693\ : InMux
    port map (
            O => \N__54081\,
            I => \N__54075\
        );

    \I__12692\ : Span4Mux_h
    port map (
            O => \N__54078\,
            I => \N__54072\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__54075\,
            I => \N__54069\
        );

    \I__12690\ : Sp12to4
    port map (
            O => \N__54072\,
            I => \N__54060\
        );

    \I__12689\ : Sp12to4
    port map (
            O => \N__54069\,
            I => \N__54060\
        );

    \I__12688\ : InMux
    port map (
            O => \N__54068\,
            I => \N__54057\
        );

    \I__12687\ : InMux
    port map (
            O => \N__54067\,
            I => \N__54052\
        );

    \I__12686\ : InMux
    port map (
            O => \N__54066\,
            I => \N__54052\
        );

    \I__12685\ : InMux
    port map (
            O => \N__54065\,
            I => \N__54049\
        );

    \I__12684\ : Span12Mux_v
    port map (
            O => \N__54060\,
            I => \N__54044\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__54057\,
            I => \N__54044\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__54052\,
            I => n21895
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__54049\,
            I => n21895
        );

    \I__12680\ : Odrv12
    port map (
            O => \N__54044\,
            I => n21895
        );

    \I__12679\ : InMux
    port map (
            O => \N__54037\,
            I => \N__54034\
        );

    \I__12678\ : LocalMux
    port map (
            O => \N__54034\,
            I => \N__54031\
        );

    \I__12677\ : Span12Mux_v
    port map (
            O => \N__54031\,
            I => \N__54028\
        );

    \I__12676\ : Odrv12
    port map (
            O => \N__54028\,
            I => buf_data_vac_8
        );

    \I__12675\ : InMux
    port map (
            O => \N__54025\,
            I => \N__54017\
        );

    \I__12674\ : InMux
    port map (
            O => \N__54024\,
            I => \N__54012\
        );

    \I__12673\ : InMux
    port map (
            O => \N__54023\,
            I => \N__54009\
        );

    \I__12672\ : InMux
    port map (
            O => \N__54022\,
            I => \N__54006\
        );

    \I__12671\ : InMux
    port map (
            O => \N__54021\,
            I => \N__54003\
        );

    \I__12670\ : InMux
    port map (
            O => \N__54020\,
            I => \N__54000\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__54017\,
            I => \N__53997\
        );

    \I__12668\ : InMux
    port map (
            O => \N__54016\,
            I => \N__53994\
        );

    \I__12667\ : InMux
    port map (
            O => \N__54015\,
            I => \N__53991\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__54012\,
            I => \N__53987\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__54009\,
            I => \N__53984\
        );

    \I__12664\ : LocalMux
    port map (
            O => \N__54006\,
            I => \N__53979\
        );

    \I__12663\ : LocalMux
    port map (
            O => \N__54003\,
            I => \N__53979\
        );

    \I__12662\ : LocalMux
    port map (
            O => \N__54000\,
            I => \N__53970\
        );

    \I__12661\ : Span4Mux_h
    port map (
            O => \N__53997\,
            I => \N__53970\
        );

    \I__12660\ : LocalMux
    port map (
            O => \N__53994\,
            I => \N__53970\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__53991\,
            I => \N__53970\
        );

    \I__12658\ : InMux
    port map (
            O => \N__53990\,
            I => \N__53967\
        );

    \I__12657\ : Span4Mux_v
    port map (
            O => \N__53987\,
            I => \N__53964\
        );

    \I__12656\ : Span4Mux_v
    port map (
            O => \N__53984\,
            I => \N__53961\
        );

    \I__12655\ : Span4Mux_v
    port map (
            O => \N__53979\,
            I => \N__53958\
        );

    \I__12654\ : Span4Mux_v
    port map (
            O => \N__53970\,
            I => \N__53953\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__53967\,
            I => \N__53953\
        );

    \I__12652\ : Span4Mux_h
    port map (
            O => \N__53964\,
            I => \N__53948\
        );

    \I__12651\ : Span4Mux_v
    port map (
            O => \N__53961\,
            I => \N__53948\
        );

    \I__12650\ : Span4Mux_v
    port map (
            O => \N__53958\,
            I => \N__53943\
        );

    \I__12649\ : Span4Mux_v
    port map (
            O => \N__53953\,
            I => \N__53943\
        );

    \I__12648\ : Odrv4
    port map (
            O => \N__53948\,
            I => comm_rx_buf_0
        );

    \I__12647\ : Odrv4
    port map (
            O => \N__53943\,
            I => comm_rx_buf_0
        );

    \I__12646\ : InMux
    port map (
            O => \N__53938\,
            I => \N__53935\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__53935\,
            I => \N__53932\
        );

    \I__12644\ : Span4Mux_v
    port map (
            O => \N__53932\,
            I => \N__53929\
        );

    \I__12643\ : Span4Mux_h
    port map (
            O => \N__53929\,
            I => \N__53926\
        );

    \I__12642\ : Span4Mux_v
    port map (
            O => \N__53926\,
            I => \N__53923\
        );

    \I__12641\ : Odrv4
    port map (
            O => \N__53923\,
            I => comm_buf_4_0
        );

    \I__12640\ : InMux
    port map (
            O => \N__53920\,
            I => \N__53917\
        );

    \I__12639\ : LocalMux
    port map (
            O => \N__53917\,
            I => \N__53914\
        );

    \I__12638\ : Span4Mux_v
    port map (
            O => \N__53914\,
            I => \N__53911\
        );

    \I__12637\ : Odrv4
    port map (
            O => \N__53911\,
            I => buf_data_vac_15
        );

    \I__12636\ : InMux
    port map (
            O => \N__53908\,
            I => \N__53905\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53902\
        );

    \I__12634\ : Span12Mux_v
    port map (
            O => \N__53902\,
            I => \N__53899\
        );

    \I__12633\ : Odrv12
    port map (
            O => \N__53899\,
            I => comm_buf_4_7
        );

    \I__12632\ : InMux
    port map (
            O => \N__53896\,
            I => \N__53890\
        );

    \I__12631\ : InMux
    port map (
            O => \N__53895\,
            I => \N__53887\
        );

    \I__12630\ : CascadeMux
    port map (
            O => \N__53894\,
            I => \N__53884\
        );

    \I__12629\ : CascadeMux
    port map (
            O => \N__53893\,
            I => \N__53880\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__53890\,
            I => \N__53874\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__53887\,
            I => \N__53874\
        );

    \I__12626\ : InMux
    port map (
            O => \N__53884\,
            I => \N__53871\
        );

    \I__12625\ : InMux
    port map (
            O => \N__53883\,
            I => \N__53868\
        );

    \I__12624\ : InMux
    port map (
            O => \N__53880\,
            I => \N__53865\
        );

    \I__12623\ : InMux
    port map (
            O => \N__53879\,
            I => \N__53862\
        );

    \I__12622\ : Span4Mux_v
    port map (
            O => \N__53874\,
            I => \N__53857\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__53871\,
            I => \N__53857\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__53868\,
            I => \N__53852\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__53865\,
            I => \N__53847\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__53862\,
            I => \N__53847\
        );

    \I__12617\ : Span4Mux_h
    port map (
            O => \N__53857\,
            I => \N__53844\
        );

    \I__12616\ : InMux
    port map (
            O => \N__53856\,
            I => \N__53841\
        );

    \I__12615\ : InMux
    port map (
            O => \N__53855\,
            I => \N__53838\
        );

    \I__12614\ : Span4Mux_v
    port map (
            O => \N__53852\,
            I => \N__53834\
        );

    \I__12613\ : Span12Mux_v
    port map (
            O => \N__53847\,
            I => \N__53827\
        );

    \I__12612\ : Sp12to4
    port map (
            O => \N__53844\,
            I => \N__53827\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__53841\,
            I => \N__53827\
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__53838\,
            I => \N__53824\
        );

    \I__12609\ : InMux
    port map (
            O => \N__53837\,
            I => \N__53821\
        );

    \I__12608\ : Odrv4
    port map (
            O => \N__53834\,
            I => comm_rx_buf_6
        );

    \I__12607\ : Odrv12
    port map (
            O => \N__53827\,
            I => comm_rx_buf_6
        );

    \I__12606\ : Odrv12
    port map (
            O => \N__53824\,
            I => comm_rx_buf_6
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__53821\,
            I => comm_rx_buf_6
        );

    \I__12604\ : InMux
    port map (
            O => \N__53812\,
            I => \N__53809\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__53809\,
            I => \N__53806\
        );

    \I__12602\ : Span4Mux_h
    port map (
            O => \N__53806\,
            I => \N__53803\
        );

    \I__12601\ : Odrv4
    port map (
            O => \N__53803\,
            I => buf_data_vac_14
        );

    \I__12600\ : InMux
    port map (
            O => \N__53800\,
            I => \N__53797\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__53797\,
            I => \N__53794\
        );

    \I__12598\ : Span4Mux_v
    port map (
            O => \N__53794\,
            I => \N__53791\
        );

    \I__12597\ : Sp12to4
    port map (
            O => \N__53791\,
            I => \N__53788\
        );

    \I__12596\ : Odrv12
    port map (
            O => \N__53788\,
            I => comm_buf_4_6
        );

    \I__12595\ : InMux
    port map (
            O => \N__53785\,
            I => \N__53782\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__53782\,
            I => \N__53772\
        );

    \I__12593\ : InMux
    port map (
            O => \N__53781\,
            I => \N__53756\
        );

    \I__12592\ : InMux
    port map (
            O => \N__53780\,
            I => \N__53756\
        );

    \I__12591\ : InMux
    port map (
            O => \N__53779\,
            I => \N__53756\
        );

    \I__12590\ : InMux
    port map (
            O => \N__53778\,
            I => \N__53756\
        );

    \I__12589\ : InMux
    port map (
            O => \N__53777\,
            I => \N__53756\
        );

    \I__12588\ : InMux
    port map (
            O => \N__53776\,
            I => \N__53756\
        );

    \I__12587\ : InMux
    port map (
            O => \N__53775\,
            I => \N__53756\
        );

    \I__12586\ : Span4Mux_v
    port map (
            O => \N__53772\,
            I => \N__53753\
        );

    \I__12585\ : InMux
    port map (
            O => \N__53771\,
            I => \N__53750\
        );

    \I__12584\ : LocalMux
    port map (
            O => \N__53756\,
            I => \N__53747\
        );

    \I__12583\ : Odrv4
    port map (
            O => \N__53753\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__53750\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__12581\ : Odrv12
    port map (
            O => \N__53747\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__12580\ : InMux
    port map (
            O => \N__53740\,
            I => \N__53730\
        );

    \I__12579\ : InMux
    port map (
            O => \N__53739\,
            I => \N__53715\
        );

    \I__12578\ : InMux
    port map (
            O => \N__53738\,
            I => \N__53715\
        );

    \I__12577\ : InMux
    port map (
            O => \N__53737\,
            I => \N__53715\
        );

    \I__12576\ : InMux
    port map (
            O => \N__53736\,
            I => \N__53715\
        );

    \I__12575\ : InMux
    port map (
            O => \N__53735\,
            I => \N__53715\
        );

    \I__12574\ : InMux
    port map (
            O => \N__53734\,
            I => \N__53715\
        );

    \I__12573\ : InMux
    port map (
            O => \N__53733\,
            I => \N__53715\
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__53730\,
            I => \comm_spi.n18536\
        );

    \I__12571\ : LocalMux
    port map (
            O => \N__53715\,
            I => \comm_spi.n18536\
        );

    \I__12570\ : ClkMux
    port map (
            O => \N__53710\,
            I => \N__53707\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__53707\,
            I => \N__53703\
        );

    \I__12568\ : ClkMux
    port map (
            O => \N__53706\,
            I => \N__53700\
        );

    \I__12567\ : Span4Mux_h
    port map (
            O => \N__53703\,
            I => \N__53692\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__53700\,
            I => \N__53692\
        );

    \I__12565\ : ClkMux
    port map (
            O => \N__53699\,
            I => \N__53685\
        );

    \I__12564\ : ClkMux
    port map (
            O => \N__53698\,
            I => \N__53682\
        );

    \I__12563\ : ClkMux
    port map (
            O => \N__53697\,
            I => \N__53679\
        );

    \I__12562\ : Span4Mux_v
    port map (
            O => \N__53692\,
            I => \N__53674\
        );

    \I__12561\ : ClkMux
    port map (
            O => \N__53691\,
            I => \N__53671\
        );

    \I__12560\ : ClkMux
    port map (
            O => \N__53690\,
            I => \N__53667\
        );

    \I__12559\ : ClkMux
    port map (
            O => \N__53689\,
            I => \N__53662\
        );

    \I__12558\ : ClkMux
    port map (
            O => \N__53688\,
            I => \N__53659\
        );

    \I__12557\ : LocalMux
    port map (
            O => \N__53685\,
            I => \N__53656\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__53682\,
            I => \N__53653\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__53679\,
            I => \N__53650\
        );

    \I__12554\ : ClkMux
    port map (
            O => \N__53678\,
            I => \N__53647\
        );

    \I__12553\ : ClkMux
    port map (
            O => \N__53677\,
            I => \N__53644\
        );

    \I__12552\ : Span4Mux_h
    port map (
            O => \N__53674\,
            I => \N__53639\
        );

    \I__12551\ : LocalMux
    port map (
            O => \N__53671\,
            I => \N__53639\
        );

    \I__12550\ : ClkMux
    port map (
            O => \N__53670\,
            I => \N__53635\
        );

    \I__12549\ : LocalMux
    port map (
            O => \N__53667\,
            I => \N__53631\
        );

    \I__12548\ : ClkMux
    port map (
            O => \N__53666\,
            I => \N__53628\
        );

    \I__12547\ : ClkMux
    port map (
            O => \N__53665\,
            I => \N__53624\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__53662\,
            I => \N__53621\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__53659\,
            I => \N__53618\
        );

    \I__12544\ : Span4Mux_v
    port map (
            O => \N__53656\,
            I => \N__53614\
        );

    \I__12543\ : Span4Mux_v
    port map (
            O => \N__53653\,
            I => \N__53609\
        );

    \I__12542\ : Span4Mux_v
    port map (
            O => \N__53650\,
            I => \N__53609\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__53647\,
            I => \N__53606\
        );

    \I__12540\ : LocalMux
    port map (
            O => \N__53644\,
            I => \N__53603\
        );

    \I__12539\ : Span4Mux_v
    port map (
            O => \N__53639\,
            I => \N__53598\
        );

    \I__12538\ : ClkMux
    port map (
            O => \N__53638\,
            I => \N__53595\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__53635\,
            I => \N__53592\
        );

    \I__12536\ : ClkMux
    port map (
            O => \N__53634\,
            I => \N__53589\
        );

    \I__12535\ : Span4Mux_h
    port map (
            O => \N__53631\,
            I => \N__53583\
        );

    \I__12534\ : LocalMux
    port map (
            O => \N__53628\,
            I => \N__53583\
        );

    \I__12533\ : ClkMux
    port map (
            O => \N__53627\,
            I => \N__53580\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__53624\,
            I => \N__53577\
        );

    \I__12531\ : Span4Mux_h
    port map (
            O => \N__53621\,
            I => \N__53572\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__53618\,
            I => \N__53572\
        );

    \I__12529\ : ClkMux
    port map (
            O => \N__53617\,
            I => \N__53569\
        );

    \I__12528\ : Span4Mux_h
    port map (
            O => \N__53614\,
            I => \N__53561\
        );

    \I__12527\ : Span4Mux_v
    port map (
            O => \N__53609\,
            I => \N__53561\
        );

    \I__12526\ : Span4Mux_v
    port map (
            O => \N__53606\,
            I => \N__53561\
        );

    \I__12525\ : Span4Mux_v
    port map (
            O => \N__53603\,
            I => \N__53558\
        );

    \I__12524\ : ClkMux
    port map (
            O => \N__53602\,
            I => \N__53555\
        );

    \I__12523\ : ClkMux
    port map (
            O => \N__53601\,
            I => \N__53552\
        );

    \I__12522\ : Span4Mux_v
    port map (
            O => \N__53598\,
            I => \N__53547\
        );

    \I__12521\ : LocalMux
    port map (
            O => \N__53595\,
            I => \N__53547\
        );

    \I__12520\ : Span4Mux_v
    port map (
            O => \N__53592\,
            I => \N__53542\
        );

    \I__12519\ : LocalMux
    port map (
            O => \N__53589\,
            I => \N__53542\
        );

    \I__12518\ : ClkMux
    port map (
            O => \N__53588\,
            I => \N__53539\
        );

    \I__12517\ : Span4Mux_v
    port map (
            O => \N__53583\,
            I => \N__53534\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__53580\,
            I => \N__53534\
        );

    \I__12515\ : Span4Mux_h
    port map (
            O => \N__53577\,
            I => \N__53531\
        );

    \I__12514\ : Span4Mux_h
    port map (
            O => \N__53572\,
            I => \N__53526\
        );

    \I__12513\ : LocalMux
    port map (
            O => \N__53569\,
            I => \N__53526\
        );

    \I__12512\ : ClkMux
    port map (
            O => \N__53568\,
            I => \N__53523\
        );

    \I__12511\ : Span4Mux_h
    port map (
            O => \N__53561\,
            I => \N__53520\
        );

    \I__12510\ : Span4Mux_v
    port map (
            O => \N__53558\,
            I => \N__53517\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__53555\,
            I => \N__53514\
        );

    \I__12508\ : LocalMux
    port map (
            O => \N__53552\,
            I => \N__53511\
        );

    \I__12507\ : Span4Mux_v
    port map (
            O => \N__53547\,
            I => \N__53504\
        );

    \I__12506\ : Span4Mux_h
    port map (
            O => \N__53542\,
            I => \N__53504\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__53539\,
            I => \N__53504\
        );

    \I__12504\ : Span4Mux_h
    port map (
            O => \N__53534\,
            I => \N__53501\
        );

    \I__12503\ : Span4Mux_h
    port map (
            O => \N__53531\,
            I => \N__53496\
        );

    \I__12502\ : Span4Mux_v
    port map (
            O => \N__53526\,
            I => \N__53496\
        );

    \I__12501\ : LocalMux
    port map (
            O => \N__53523\,
            I => \N__53493\
        );

    \I__12500\ : Span4Mux_v
    port map (
            O => \N__53520\,
            I => \N__53490\
        );

    \I__12499\ : Span4Mux_h
    port map (
            O => \N__53517\,
            I => \N__53485\
        );

    \I__12498\ : Span4Mux_v
    port map (
            O => \N__53514\,
            I => \N__53485\
        );

    \I__12497\ : Span4Mux_v
    port map (
            O => \N__53511\,
            I => \N__53480\
        );

    \I__12496\ : Span4Mux_h
    port map (
            O => \N__53504\,
            I => \N__53480\
        );

    \I__12495\ : Sp12to4
    port map (
            O => \N__53501\,
            I => \N__53473\
        );

    \I__12494\ : Sp12to4
    port map (
            O => \N__53496\,
            I => \N__53473\
        );

    \I__12493\ : Sp12to4
    port map (
            O => \N__53493\,
            I => \N__53473\
        );

    \I__12492\ : Odrv4
    port map (
            O => \N__53490\,
            I => \comm_spi.iclk\
        );

    \I__12491\ : Odrv4
    port map (
            O => \N__53485\,
            I => \comm_spi.iclk\
        );

    \I__12490\ : Odrv4
    port map (
            O => \N__53480\,
            I => \comm_spi.iclk\
        );

    \I__12489\ : Odrv12
    port map (
            O => \N__53473\,
            I => \comm_spi.iclk\
        );

    \I__12488\ : InMux
    port map (
            O => \N__53464\,
            I => \N__53461\
        );

    \I__12487\ : LocalMux
    port map (
            O => \N__53461\,
            I => \N__53458\
        );

    \I__12486\ : Odrv4
    port map (
            O => \N__53458\,
            I => n22330
        );

    \I__12485\ : CascadeMux
    port map (
            O => \N__53455\,
            I => \N__53452\
        );

    \I__12484\ : InMux
    port map (
            O => \N__53452\,
            I => \N__53449\
        );

    \I__12483\ : LocalMux
    port map (
            O => \N__53449\,
            I => n22329
        );

    \I__12482\ : InMux
    port map (
            O => \N__53446\,
            I => \N__53443\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__53443\,
            I => \N__53440\
        );

    \I__12480\ : Span4Mux_v
    port map (
            O => \N__53440\,
            I => \N__53435\
        );

    \I__12479\ : InMux
    port map (
            O => \N__53439\,
            I => \N__53432\
        );

    \I__12478\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53429\
        );

    \I__12477\ : Span4Mux_h
    port map (
            O => \N__53435\,
            I => \N__53426\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__53432\,
            I => n15261
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__53429\,
            I => n15261
        );

    \I__12474\ : Odrv4
    port map (
            O => \N__53426\,
            I => n15261
        );

    \I__12473\ : CascadeMux
    port map (
            O => \N__53419\,
            I => \n22321_cascade_\
        );

    \I__12472\ : CascadeMux
    port map (
            O => \N__53416\,
            I => \N__53413\
        );

    \I__12471\ : InMux
    port map (
            O => \N__53413\,
            I => \N__53410\
        );

    \I__12470\ : LocalMux
    port map (
            O => \N__53410\,
            I => \N__53406\
        );

    \I__12469\ : InMux
    port map (
            O => \N__53409\,
            I => \N__53403\
        );

    \I__12468\ : Odrv4
    port map (
            O => \N__53406\,
            I => n14851
        );

    \I__12467\ : LocalMux
    port map (
            O => \N__53403\,
            I => n14851
        );

    \I__12466\ : InMux
    port map (
            O => \N__53398\,
            I => \N__53395\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__53395\,
            I => n22352
        );

    \I__12464\ : InMux
    port map (
            O => \N__53392\,
            I => \N__53388\
        );

    \I__12463\ : InMux
    port map (
            O => \N__53391\,
            I => \N__53385\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__53388\,
            I => dds0_mclkcnt_6
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__53385\,
            I => dds0_mclkcnt_6
        );

    \I__12460\ : IoInMux
    port map (
            O => \N__53380\,
            I => \N__53377\
        );

    \I__12459\ : LocalMux
    port map (
            O => \N__53377\,
            I => \N__53374\
        );

    \I__12458\ : Span4Mux_s3_v
    port map (
            O => \N__53374\,
            I => \N__53371\
        );

    \I__12457\ : Span4Mux_v
    port map (
            O => \N__53371\,
            I => \N__53368\
        );

    \I__12456\ : Sp12to4
    port map (
            O => \N__53368\,
            I => \N__53365\
        );

    \I__12455\ : Span12Mux_v
    port map (
            O => \N__53365\,
            I => \N__53361\
        );

    \I__12454\ : InMux
    port map (
            O => \N__53364\,
            I => \N__53358\
        );

    \I__12453\ : Odrv12
    port map (
            O => \N__53361\,
            I => \DDS_MCLK\
        );

    \I__12452\ : LocalMux
    port map (
            O => \N__53358\,
            I => \DDS_MCLK\
        );

    \I__12451\ : CascadeMux
    port map (
            O => \N__53353\,
            I => \n6888_cascade_\
        );

    \I__12450\ : InMux
    port map (
            O => \N__53350\,
            I => \N__53346\
        );

    \I__12449\ : InMux
    port map (
            O => \N__53349\,
            I => \N__53343\
        );

    \I__12448\ : LocalMux
    port map (
            O => \N__53346\,
            I => n21865
        );

    \I__12447\ : LocalMux
    port map (
            O => \N__53343\,
            I => n21865
        );

    \I__12446\ : CascadeMux
    port map (
            O => \N__53338\,
            I => \N__53335\
        );

    \I__12445\ : InMux
    port map (
            O => \N__53335\,
            I => \N__53332\
        );

    \I__12444\ : LocalMux
    port map (
            O => \N__53332\,
            I => \N__53329\
        );

    \I__12443\ : Odrv4
    port map (
            O => \N__53329\,
            I => n21981
        );

    \I__12442\ : InMux
    port map (
            O => \N__53326\,
            I => \N__53323\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__53323\,
            I => n22027
        );

    \I__12440\ : InMux
    port map (
            O => \N__53320\,
            I => \N__53317\
        );

    \I__12439\ : LocalMux
    port map (
            O => \N__53317\,
            I => n22018
        );

    \I__12438\ : InMux
    port map (
            O => \N__53314\,
            I => \N__53310\
        );

    \I__12437\ : InMux
    port map (
            O => \N__53313\,
            I => \N__53307\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__53310\,
            I => dds0_mclkcnt_3
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__53307\,
            I => dds0_mclkcnt_3
        );

    \I__12434\ : InMux
    port map (
            O => \N__53302\,
            I => \N__53298\
        );

    \I__12433\ : InMux
    port map (
            O => \N__53301\,
            I => \N__53295\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__53298\,
            I => dds0_mclkcnt_5
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__53295\,
            I => dds0_mclkcnt_5
        );

    \I__12430\ : CascadeMux
    port map (
            O => \N__53290\,
            I => \N__53287\
        );

    \I__12429\ : InMux
    port map (
            O => \N__53287\,
            I => \N__53283\
        );

    \I__12428\ : InMux
    port map (
            O => \N__53286\,
            I => \N__53280\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__53283\,
            I => \N__53277\
        );

    \I__12426\ : LocalMux
    port map (
            O => \N__53280\,
            I => dds0_mclkcnt_1
        );

    \I__12425\ : Odrv4
    port map (
            O => \N__53277\,
            I => dds0_mclkcnt_1
        );

    \I__12424\ : InMux
    port map (
            O => \N__53272\,
            I => \N__53268\
        );

    \I__12423\ : InMux
    port map (
            O => \N__53271\,
            I => \N__53265\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__53268\,
            I => dds0_mclkcnt_4
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__53265\,
            I => dds0_mclkcnt_4
        );

    \I__12420\ : InMux
    port map (
            O => \N__53260\,
            I => \N__53256\
        );

    \I__12419\ : InMux
    port map (
            O => \N__53259\,
            I => \N__53253\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__53256\,
            I => \N__53250\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__53253\,
            I => dds0_mclkcnt_7
        );

    \I__12416\ : Odrv4
    port map (
            O => \N__53250\,
            I => dds0_mclkcnt_7
        );

    \I__12415\ : InMux
    port map (
            O => \N__53245\,
            I => \N__53241\
        );

    \I__12414\ : InMux
    port map (
            O => \N__53244\,
            I => \N__53238\
        );

    \I__12413\ : LocalMux
    port map (
            O => \N__53241\,
            I => dds0_mclkcnt_0
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__53238\,
            I => dds0_mclkcnt_0
        );

    \I__12411\ : CascadeMux
    port map (
            O => \N__53233\,
            I => \n12_adj_1685_cascade_\
        );

    \I__12410\ : InMux
    port map (
            O => \N__53230\,
            I => \N__53226\
        );

    \I__12409\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53223\
        );

    \I__12408\ : LocalMux
    port map (
            O => \N__53226\,
            I => dds0_mclkcnt_2
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__53223\,
            I => dds0_mclkcnt_2
        );

    \I__12406\ : InMux
    port map (
            O => \N__53218\,
            I => \N__53212\
        );

    \I__12405\ : InMux
    port map (
            O => \N__53217\,
            I => \N__53212\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__53212\,
            I => n21857
        );

    \I__12403\ : InMux
    port map (
            O => \N__53209\,
            I => \bfn_19_7_0_\
        );

    \I__12402\ : InMux
    port map (
            O => \N__53206\,
            I => n20819
        );

    \I__12401\ : InMux
    port map (
            O => \N__53203\,
            I => n20820
        );

    \I__12400\ : InMux
    port map (
            O => \N__53200\,
            I => n20821
        );

    \I__12399\ : InMux
    port map (
            O => \N__53197\,
            I => n20822
        );

    \I__12398\ : InMux
    port map (
            O => \N__53194\,
            I => n20823
        );

    \I__12397\ : InMux
    port map (
            O => \N__53191\,
            I => n20824
        );

    \I__12396\ : InMux
    port map (
            O => \N__53188\,
            I => n20825
        );

    \I__12395\ : InMux
    port map (
            O => \N__53185\,
            I => \N__53182\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__53182\,
            I => n10
        );

    \I__12393\ : InMux
    port map (
            O => \N__53179\,
            I => \ADC_VDC.genclk.n20757\
        );

    \I__12392\ : InMux
    port map (
            O => \N__53176\,
            I => \bfn_19_6_0_\
        );

    \I__12391\ : InMux
    port map (
            O => \N__53173\,
            I => \ADC_VDC.genclk.n20759\
        );

    \I__12390\ : InMux
    port map (
            O => \N__53170\,
            I => \ADC_VDC.genclk.n20760\
        );

    \I__12389\ : InMux
    port map (
            O => \N__53167\,
            I => \ADC_VDC.genclk.n20761\
        );

    \I__12388\ : InMux
    port map (
            O => \N__53164\,
            I => \ADC_VDC.genclk.n20762\
        );

    \I__12387\ : InMux
    port map (
            O => \N__53161\,
            I => \ADC_VDC.genclk.n20763\
        );

    \I__12386\ : InMux
    port map (
            O => \N__53158\,
            I => \ADC_VDC.genclk.n20764\
        );

    \I__12385\ : InMux
    port map (
            O => \N__53155\,
            I => \ADC_VDC.genclk.n20765\
        );

    \I__12384\ : InMux
    port map (
            O => \N__53152\,
            I => \N__53148\
        );

    \I__12383\ : InMux
    port map (
            O => \N__53151\,
            I => \N__53145\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__53148\,
            I => \N__53142\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__53145\,
            I => \N__53139\
        );

    \I__12380\ : Span4Mux_v
    port map (
            O => \N__53142\,
            I => \N__53136\
        );

    \I__12379\ : Span4Mux_h
    port map (
            O => \N__53139\,
            I => \N__53133\
        );

    \I__12378\ : Span4Mux_h
    port map (
            O => \N__53136\,
            I => \N__53130\
        );

    \I__12377\ : Span4Mux_v
    port map (
            O => \N__53133\,
            I => \N__53127\
        );

    \I__12376\ : Odrv4
    port map (
            O => \N__53130\,
            I => n7
        );

    \I__12375\ : Odrv4
    port map (
            O => \N__53127\,
            I => n7
        );

    \I__12374\ : CascadeMux
    port map (
            O => \N__53122\,
            I => \N__53119\
        );

    \I__12373\ : CascadeBuf
    port map (
            O => \N__53119\,
            I => \N__53116\
        );

    \I__12372\ : CascadeMux
    port map (
            O => \N__53116\,
            I => \N__53113\
        );

    \I__12371\ : CascadeBuf
    port map (
            O => \N__53113\,
            I => \N__53110\
        );

    \I__12370\ : CascadeMux
    port map (
            O => \N__53110\,
            I => \N__53107\
        );

    \I__12369\ : CascadeBuf
    port map (
            O => \N__53107\,
            I => \N__53104\
        );

    \I__12368\ : CascadeMux
    port map (
            O => \N__53104\,
            I => \N__53101\
        );

    \I__12367\ : CascadeBuf
    port map (
            O => \N__53101\,
            I => \N__53098\
        );

    \I__12366\ : CascadeMux
    port map (
            O => \N__53098\,
            I => \N__53095\
        );

    \I__12365\ : CascadeBuf
    port map (
            O => \N__53095\,
            I => \N__53092\
        );

    \I__12364\ : CascadeMux
    port map (
            O => \N__53092\,
            I => \N__53089\
        );

    \I__12363\ : CascadeBuf
    port map (
            O => \N__53089\,
            I => \N__53086\
        );

    \I__12362\ : CascadeMux
    port map (
            O => \N__53086\,
            I => \N__53083\
        );

    \I__12361\ : CascadeBuf
    port map (
            O => \N__53083\,
            I => \N__53079\
        );

    \I__12360\ : CascadeMux
    port map (
            O => \N__53082\,
            I => \N__53076\
        );

    \I__12359\ : CascadeMux
    port map (
            O => \N__53079\,
            I => \N__53073\
        );

    \I__12358\ : CascadeBuf
    port map (
            O => \N__53076\,
            I => \N__53070\
        );

    \I__12357\ : CascadeBuf
    port map (
            O => \N__53073\,
            I => \N__53067\
        );

    \I__12356\ : CascadeMux
    port map (
            O => \N__53070\,
            I => \N__53064\
        );

    \I__12355\ : CascadeMux
    port map (
            O => \N__53067\,
            I => \N__53061\
        );

    \I__12354\ : InMux
    port map (
            O => \N__53064\,
            I => \N__53058\
        );

    \I__12353\ : CascadeBuf
    port map (
            O => \N__53061\,
            I => \N__53055\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__53058\,
            I => \N__53052\
        );

    \I__12351\ : CascadeMux
    port map (
            O => \N__53055\,
            I => \N__53049\
        );

    \I__12350\ : Span12Mux_h
    port map (
            O => \N__53052\,
            I => \N__53046\
        );

    \I__12349\ : InMux
    port map (
            O => \N__53049\,
            I => \N__53043\
        );

    \I__12348\ : Span12Mux_v
    port map (
            O => \N__53046\,
            I => \N__53038\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__53043\,
            I => \N__53038\
        );

    \I__12346\ : Odrv12
    port map (
            O => \N__53038\,
            I => \data_index_9_N_236_0\
        );

    \I__12345\ : InMux
    port map (
            O => \N__53035\,
            I => \N__53032\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__53032\,
            I => \N__53029\
        );

    \I__12343\ : Odrv4
    port map (
            O => \N__53029\,
            I => buf_data_iac_20
        );

    \I__12342\ : InMux
    port map (
            O => \N__53026\,
            I => \N__53023\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__53023\,
            I => \N__53020\
        );

    \I__12340\ : Span12Mux_v
    port map (
            O => \N__53020\,
            I => \N__53017\
        );

    \I__12339\ : Odrv12
    port map (
            O => \N__53017\,
            I => n22500
        );

    \I__12338\ : InMux
    port map (
            O => \N__53014\,
            I => \bfn_19_5_0_\
        );

    \I__12337\ : InMux
    port map (
            O => \N__53011\,
            I => \ADC_VDC.genclk.n20751\
        );

    \I__12336\ : InMux
    port map (
            O => \N__53008\,
            I => \ADC_VDC.genclk.n20752\
        );

    \I__12335\ : InMux
    port map (
            O => \N__53005\,
            I => \ADC_VDC.genclk.n20753\
        );

    \I__12334\ : InMux
    port map (
            O => \N__53002\,
            I => \ADC_VDC.genclk.n20754\
        );

    \I__12333\ : InMux
    port map (
            O => \N__52999\,
            I => \ADC_VDC.genclk.n20755\
        );

    \I__12332\ : InMux
    port map (
            O => \N__52996\,
            I => \ADC_VDC.genclk.n20756\
        );

    \I__12331\ : CascadeMux
    port map (
            O => \N__52993\,
            I => \n22152_cascade_\
        );

    \I__12330\ : InMux
    port map (
            O => \N__52990\,
            I => \N__52987\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__52987\,
            I => \N__52984\
        );

    \I__12328\ : Sp12to4
    port map (
            O => \N__52984\,
            I => \N__52981\
        );

    \I__12327\ : Span12Mux_v
    port map (
            O => \N__52981\,
            I => \N__52978\
        );

    \I__12326\ : Span12Mux_h
    port map (
            O => \N__52978\,
            I => \N__52975\
        );

    \I__12325\ : Odrv12
    port map (
            O => \N__52975\,
            I => n22149
        );

    \I__12324\ : CascadeMux
    port map (
            O => \N__52972\,
            I => \n23444_cascade_\
        );

    \I__12323\ : InMux
    port map (
            O => \N__52969\,
            I => \N__52966\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__52966\,
            I => \N__52963\
        );

    \I__12321\ : Span4Mux_h
    port map (
            O => \N__52963\,
            I => \N__52960\
        );

    \I__12320\ : Odrv4
    port map (
            O => \N__52960\,
            I => n22148
        );

    \I__12319\ : InMux
    port map (
            O => \N__52957\,
            I => \N__52954\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__52954\,
            I => \N__52951\
        );

    \I__12317\ : Span4Mux_h
    port map (
            O => \N__52951\,
            I => \N__52948\
        );

    \I__12316\ : Span4Mux_h
    port map (
            O => \N__52948\,
            I => \N__52945\
        );

    \I__12315\ : Odrv4
    port map (
            O => \N__52945\,
            I => n111_adj_1750
        );

    \I__12314\ : CascadeMux
    port map (
            O => \N__52942\,
            I => \n23447_cascade_\
        );

    \I__12313\ : CascadeMux
    port map (
            O => \N__52939\,
            I => \comm_buf_1_7_N_559_2_cascade_\
        );

    \I__12312\ : InMux
    port map (
            O => \N__52936\,
            I => \N__52931\
        );

    \I__12311\ : CascadeMux
    port map (
            O => \N__52935\,
            I => \N__52928\
        );

    \I__12310\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52922\
        );

    \I__12309\ : LocalMux
    port map (
            O => \N__52931\,
            I => \N__52919\
        );

    \I__12308\ : InMux
    port map (
            O => \N__52928\,
            I => \N__52916\
        );

    \I__12307\ : InMux
    port map (
            O => \N__52927\,
            I => \N__52913\
        );

    \I__12306\ : InMux
    port map (
            O => \N__52926\,
            I => \N__52910\
        );

    \I__12305\ : CascadeMux
    port map (
            O => \N__52925\,
            I => \N__52906\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__52922\,
            I => \N__52901\
        );

    \I__12303\ : Span4Mux_v
    port map (
            O => \N__52919\,
            I => \N__52901\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__52916\,
            I => \N__52896\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__52913\,
            I => \N__52896\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__52910\,
            I => \N__52893\
        );

    \I__12299\ : InMux
    port map (
            O => \N__52909\,
            I => \N__52890\
        );

    \I__12298\ : InMux
    port map (
            O => \N__52906\,
            I => \N__52885\
        );

    \I__12297\ : Span4Mux_v
    port map (
            O => \N__52901\,
            I => \N__52880\
        );

    \I__12296\ : Span4Mux_v
    port map (
            O => \N__52896\,
            I => \N__52880\
        );

    \I__12295\ : Span4Mux_v
    port map (
            O => \N__52893\,
            I => \N__52875\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__52890\,
            I => \N__52875\
        );

    \I__12293\ : InMux
    port map (
            O => \N__52889\,
            I => \N__52870\
        );

    \I__12292\ : InMux
    port map (
            O => \N__52888\,
            I => \N__52870\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__52885\,
            I => \N__52867\
        );

    \I__12290\ : Span4Mux_h
    port map (
            O => \N__52880\,
            I => \N__52864\
        );

    \I__12289\ : Span4Mux_v
    port map (
            O => \N__52875\,
            I => \N__52859\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__52870\,
            I => \N__52859\
        );

    \I__12287\ : Span4Mux_h
    port map (
            O => \N__52867\,
            I => \N__52856\
        );

    \I__12286\ : Span4Mux_h
    port map (
            O => \N__52864\,
            I => \N__52853\
        );

    \I__12285\ : Span4Mux_h
    port map (
            O => \N__52859\,
            I => \N__52850\
        );

    \I__12284\ : Odrv4
    port map (
            O => \N__52856\,
            I => comm_buf_1_2
        );

    \I__12283\ : Odrv4
    port map (
            O => \N__52853\,
            I => comm_buf_1_2
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__52850\,
            I => comm_buf_1_2
        );

    \I__12281\ : InMux
    port map (
            O => \N__52843\,
            I => \N__52839\
        );

    \I__12280\ : CascadeMux
    port map (
            O => \N__52842\,
            I => \N__52836\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__52839\,
            I => \N__52833\
        );

    \I__12278\ : InMux
    port map (
            O => \N__52836\,
            I => \N__52829\
        );

    \I__12277\ : Span4Mux_h
    port map (
            O => \N__52833\,
            I => \N__52826\
        );

    \I__12276\ : InMux
    port map (
            O => \N__52832\,
            I => \N__52823\
        );

    \I__12275\ : LocalMux
    port map (
            O => \N__52829\,
            I => req_data_cnt_2
        );

    \I__12274\ : Odrv4
    port map (
            O => \N__52826\,
            I => req_data_cnt_2
        );

    \I__12273\ : LocalMux
    port map (
            O => \N__52823\,
            I => req_data_cnt_2
        );

    \I__12272\ : CascadeMux
    port map (
            O => \N__52816\,
            I => \N__52813\
        );

    \I__12271\ : InMux
    port map (
            O => \N__52813\,
            I => \N__52808\
        );

    \I__12270\ : InMux
    port map (
            O => \N__52812\,
            I => \N__52805\
        );

    \I__12269\ : CascadeMux
    port map (
            O => \N__52811\,
            I => \N__52802\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__52808\,
            I => \N__52799\
        );

    \I__12267\ : LocalMux
    port map (
            O => \N__52805\,
            I => \N__52796\
        );

    \I__12266\ : InMux
    port map (
            O => \N__52802\,
            I => \N__52793\
        );

    \I__12265\ : Odrv4
    port map (
            O => \N__52799\,
            I => \acadc_skipCount_2\
        );

    \I__12264\ : Odrv12
    port map (
            O => \N__52796\,
            I => \acadc_skipCount_2\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__52793\,
            I => \acadc_skipCount_2\
        );

    \I__12262\ : InMux
    port map (
            O => \N__52786\,
            I => \N__52783\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__52783\,
            I => n22151
        );

    \I__12260\ : IoInMux
    port map (
            O => \N__52780\,
            I => \N__52776\
        );

    \I__12259\ : InMux
    port map (
            O => \N__52779\,
            I => \N__52773\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__52776\,
            I => \N__52770\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__52773\,
            I => \N__52767\
        );

    \I__12256\ : Span4Mux_s3_v
    port map (
            O => \N__52770\,
            I => \N__52764\
        );

    \I__12255\ : Span4Mux_h
    port map (
            O => \N__52767\,
            I => \N__52760\
        );

    \I__12254\ : Span4Mux_v
    port map (
            O => \N__52764\,
            I => \N__52757\
        );

    \I__12253\ : InMux
    port map (
            O => \N__52763\,
            I => \N__52754\
        );

    \I__12252\ : Span4Mux_h
    port map (
            O => \N__52760\,
            I => \N__52751\
        );

    \I__12251\ : Odrv4
    port map (
            O => \N__52757\,
            I => \SELIRNG1\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__52754\,
            I => \SELIRNG1\
        );

    \I__12249\ : Odrv4
    port map (
            O => \N__52751\,
            I => \SELIRNG1\
        );

    \I__12248\ : InMux
    port map (
            O => \N__52744\,
            I => \N__52739\
        );

    \I__12247\ : CascadeMux
    port map (
            O => \N__52743\,
            I => \N__52736\
        );

    \I__12246\ : InMux
    port map (
            O => \N__52742\,
            I => \N__52733\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__52739\,
            I => \N__52730\
        );

    \I__12244\ : InMux
    port map (
            O => \N__52736\,
            I => \N__52727\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__52733\,
            I => \acadc_skipCount_11\
        );

    \I__12242\ : Odrv12
    port map (
            O => \N__52730\,
            I => \acadc_skipCount_11\
        );

    \I__12241\ : LocalMux
    port map (
            O => \N__52727\,
            I => \acadc_skipCount_11\
        );

    \I__12240\ : InMux
    port map (
            O => \N__52720\,
            I => \N__52717\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__52717\,
            I => \N__52713\
        );

    \I__12238\ : InMux
    port map (
            O => \N__52716\,
            I => \N__52710\
        );

    \I__12237\ : Span4Mux_v
    port map (
            O => \N__52713\,
            I => \N__52705\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52705\
        );

    \I__12235\ : Span4Mux_h
    port map (
            O => \N__52705\,
            I => \N__52701\
        );

    \I__12234\ : InMux
    port map (
            O => \N__52704\,
            I => \N__52698\
        );

    \I__12233\ : Span4Mux_h
    port map (
            O => \N__52701\,
            I => \N__52695\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__52698\,
            I => buf_adcdata_iac_9
        );

    \I__12231\ : Odrv4
    port map (
            O => \N__52695\,
            I => buf_adcdata_iac_9
        );

    \I__12230\ : InMux
    port map (
            O => \N__52690\,
            I => \N__52687\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__52687\,
            I => \N__52684\
        );

    \I__12228\ : Odrv12
    port map (
            O => \N__52684\,
            I => n16_adj_1751
        );

    \I__12227\ : InMux
    port map (
            O => \N__52681\,
            I => \N__52678\
        );

    \I__12226\ : LocalMux
    port map (
            O => \N__52678\,
            I => \N__52675\
        );

    \I__12225\ : Span4Mux_v
    port map (
            O => \N__52675\,
            I => \N__52672\
        );

    \I__12224\ : Odrv4
    port map (
            O => \N__52672\,
            I => n22136
        );

    \I__12223\ : InMux
    port map (
            O => \N__52669\,
            I => \N__52666\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__52666\,
            I => \N__52663\
        );

    \I__12221\ : Span12Mux_h
    port map (
            O => \N__52663\,
            I => \N__52660\
        );

    \I__12220\ : Span12Mux_v
    port map (
            O => \N__52660\,
            I => \N__52655\
        );

    \I__12219\ : InMux
    port map (
            O => \N__52659\,
            I => \N__52652\
        );

    \I__12218\ : InMux
    port map (
            O => \N__52658\,
            I => \N__52649\
        );

    \I__12217\ : Odrv12
    port map (
            O => \N__52655\,
            I => wdtick_flag
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__52652\,
            I => wdtick_flag
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__52649\,
            I => wdtick_flag
        );

    \I__12214\ : CascadeMux
    port map (
            O => \N__52642\,
            I => \N__52639\
        );

    \I__12213\ : InMux
    port map (
            O => \N__52639\,
            I => \N__52635\
        );

    \I__12212\ : InMux
    port map (
            O => \N__52638\,
            I => \N__52632\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__52635\,
            I => \N__52629\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__52632\,
            I => \N__52626\
        );

    \I__12209\ : Span4Mux_h
    port map (
            O => \N__52629\,
            I => \N__52622\
        );

    \I__12208\ : Span4Mux_v
    port map (
            O => \N__52626\,
            I => \N__52619\
        );

    \I__12207\ : InMux
    port map (
            O => \N__52625\,
            I => \N__52616\
        );

    \I__12206\ : Span4Mux_h
    port map (
            O => \N__52622\,
            I => \N__52613\
        );

    \I__12205\ : Odrv4
    port map (
            O => \N__52619\,
            I => buf_control_0
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__52616\,
            I => buf_control_0
        );

    \I__12203\ : Odrv4
    port map (
            O => \N__52613\,
            I => buf_control_0
        );

    \I__12202\ : IoInMux
    port map (
            O => \N__52606\,
            I => \N__52603\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52600\
        );

    \I__12200\ : Span4Mux_s1_v
    port map (
            O => \N__52600\,
            I => \N__52597\
        );

    \I__12199\ : Span4Mux_h
    port map (
            O => \N__52597\,
            I => \N__52594\
        );

    \I__12198\ : Span4Mux_v
    port map (
            O => \N__52594\,
            I => \N__52591\
        );

    \I__12197\ : Odrv4
    port map (
            O => \N__52591\,
            I => \CONT_SD\
        );

    \I__12196\ : InMux
    port map (
            O => \N__52588\,
            I => \N__52584\
        );

    \I__12195\ : InMux
    port map (
            O => \N__52587\,
            I => \N__52581\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__52584\,
            I => \N__52578\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__52581\,
            I => \N__52575\
        );

    \I__12192\ : Span4Mux_h
    port map (
            O => \N__52578\,
            I => \N__52572\
        );

    \I__12191\ : Odrv4
    port map (
            O => \N__52575\,
            I => n8_adj_1605
        );

    \I__12190\ : Odrv4
    port map (
            O => \N__52572\,
            I => n8_adj_1605
        );

    \I__12189\ : InMux
    port map (
            O => \N__52567\,
            I => \N__52564\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__52564\,
            I => \N__52560\
        );

    \I__12187\ : InMux
    port map (
            O => \N__52563\,
            I => \N__52557\
        );

    \I__12186\ : Span4Mux_h
    port map (
            O => \N__52560\,
            I => \N__52554\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__52557\,
            I => data_idxvec_4
        );

    \I__12184\ : Odrv4
    port map (
            O => \N__52554\,
            I => data_idxvec_4
        );

    \I__12183\ : InMux
    port map (
            O => \N__52549\,
            I => \N__52546\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__52546\,
            I => \N__52542\
        );

    \I__12181\ : InMux
    port map (
            O => \N__52545\,
            I => \N__52538\
        );

    \I__12180\ : Span4Mux_h
    port map (
            O => \N__52542\,
            I => \N__52535\
        );

    \I__12179\ : InMux
    port map (
            O => \N__52541\,
            I => \N__52532\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__52538\,
            I => data_cntvec_4
        );

    \I__12177\ : Odrv4
    port map (
            O => \N__52535\,
            I => data_cntvec_4
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__52532\,
            I => data_cntvec_4
        );

    \I__12175\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52522\
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__52522\,
            I => \N__52519\
        );

    \I__12173\ : Odrv12
    port map (
            O => \N__52519\,
            I => n22301
        );

    \I__12172\ : CascadeMux
    port map (
            O => \N__52516\,
            I => \n26_adj_1735_cascade_\
        );

    \I__12171\ : CascadeMux
    port map (
            O => \N__52513\,
            I => \N__52509\
        );

    \I__12170\ : InMux
    port map (
            O => \N__52512\,
            I => \N__52506\
        );

    \I__12169\ : InMux
    port map (
            O => \N__52509\,
            I => \N__52502\
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52499\
        );

    \I__12167\ : InMux
    port map (
            O => \N__52505\,
            I => \N__52496\
        );

    \I__12166\ : LocalMux
    port map (
            O => \N__52502\,
            I => \acadc_skipCount_4\
        );

    \I__12165\ : Odrv4
    port map (
            O => \N__52499\,
            I => \acadc_skipCount_4\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__52496\,
            I => \acadc_skipCount_4\
        );

    \I__12163\ : CascadeMux
    port map (
            O => \N__52489\,
            I => \n23318_cascade_\
        );

    \I__12162\ : InMux
    port map (
            O => \N__52486\,
            I => \N__52483\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__52483\,
            I => \N__52478\
        );

    \I__12160\ : InMux
    port map (
            O => \N__52482\,
            I => \N__52475\
        );

    \I__12159\ : InMux
    port map (
            O => \N__52481\,
            I => \N__52472\
        );

    \I__12158\ : Span4Mux_v
    port map (
            O => \N__52478\,
            I => \N__52467\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__52475\,
            I => \N__52467\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__52472\,
            I => req_data_cnt_4
        );

    \I__12155\ : Odrv4
    port map (
            O => \N__52467\,
            I => req_data_cnt_4
        );

    \I__12154\ : InMux
    port map (
            O => \N__52462\,
            I => \N__52459\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__52459\,
            I => \N__52456\
        );

    \I__12152\ : Span4Mux_h
    port map (
            O => \N__52456\,
            I => \N__52453\
        );

    \I__12151\ : Span4Mux_h
    port map (
            O => \N__52453\,
            I => \N__52450\
        );

    \I__12150\ : Odrv4
    port map (
            O => \N__52450\,
            I => n23441
        );

    \I__12149\ : CascadeMux
    port map (
            O => \N__52447\,
            I => \n23321_cascade_\
        );

    \I__12148\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52441\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__52441\,
            I => \N__52438\
        );

    \I__12146\ : Span4Mux_v
    port map (
            O => \N__52438\,
            I => \N__52435\
        );

    \I__12145\ : Span4Mux_h
    port map (
            O => \N__52435\,
            I => \N__52432\
        );

    \I__12144\ : Span4Mux_h
    port map (
            O => \N__52432\,
            I => \N__52429\
        );

    \I__12143\ : Odrv4
    port map (
            O => \N__52429\,
            I => n111_adj_1737
        );

    \I__12142\ : CascadeMux
    port map (
            O => \N__52426\,
            I => \n30_adj_1736_cascade_\
        );

    \I__12141\ : CascadeMux
    port map (
            O => \N__52423\,
            I => \comm_buf_1_7_N_559_4_cascade_\
        );

    \I__12140\ : InMux
    port map (
            O => \N__52420\,
            I => \N__52416\
        );

    \I__12139\ : InMux
    port map (
            O => \N__52419\,
            I => \N__52413\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__52416\,
            I => \N__52408\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__52413\,
            I => \N__52408\
        );

    \I__12136\ : Odrv4
    port map (
            O => \N__52408\,
            I => data_idxvec_2
        );

    \I__12135\ : CascadeMux
    port map (
            O => \N__52405\,
            I => \N__52402\
        );

    \I__12134\ : InMux
    port map (
            O => \N__52402\,
            I => \N__52399\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__52399\,
            I => \N__52394\
        );

    \I__12132\ : InMux
    port map (
            O => \N__52398\,
            I => \N__52391\
        );

    \I__12131\ : InMux
    port map (
            O => \N__52397\,
            I => \N__52388\
        );

    \I__12130\ : Span4Mux_h
    port map (
            O => \N__52394\,
            I => \N__52385\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__52391\,
            I => data_cntvec_2
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__52388\,
            I => data_cntvec_2
        );

    \I__12127\ : Odrv4
    port map (
            O => \N__52385\,
            I => data_cntvec_2
        );

    \I__12126\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52375\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__52375\,
            I => \N__52372\
        );

    \I__12124\ : Span4Mux_v
    port map (
            O => \N__52372\,
            I => \N__52369\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__52369\,
            I => buf_data_iac_10
        );

    \I__12122\ : CascadeMux
    port map (
            O => \N__52366\,
            I => \n26_adj_1748_cascade_\
        );

    \I__12121\ : CascadeMux
    port map (
            O => \N__52363\,
            I => \comm_buf_1_7_N_559_5_cascade_\
        );

    \I__12120\ : InMux
    port map (
            O => \N__52360\,
            I => \N__52357\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__52357\,
            I => \N__52354\
        );

    \I__12118\ : Span4Mux_v
    port map (
            O => \N__52354\,
            I => \N__52351\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__52351\,
            I => \N__52348\
        );

    \I__12116\ : Span4Mux_h
    port map (
            O => \N__52348\,
            I => \N__52345\
        );

    \I__12115\ : Odrv4
    port map (
            O => \N__52345\,
            I => n16_adj_1728
        );

    \I__12114\ : CascadeMux
    port map (
            O => \N__52342\,
            I => \N__52338\
        );

    \I__12113\ : InMux
    port map (
            O => \N__52341\,
            I => \N__52335\
        );

    \I__12112\ : InMux
    port map (
            O => \N__52338\,
            I => \N__52332\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__52335\,
            I => \N__52329\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__52332\,
            I => \N__52326\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__52329\,
            I => \N__52323\
        );

    \I__12108\ : Span4Mux_v
    port map (
            O => \N__52326\,
            I => \N__52320\
        );

    \I__12107\ : Sp12to4
    port map (
            O => \N__52323\,
            I => \N__52316\
        );

    \I__12106\ : Span4Mux_h
    port map (
            O => \N__52320\,
            I => \N__52313\
        );

    \I__12105\ : InMux
    port map (
            O => \N__52319\,
            I => \N__52310\
        );

    \I__12104\ : Span12Mux_h
    port map (
            O => \N__52316\,
            I => \N__52307\
        );

    \I__12103\ : Span4Mux_h
    port map (
            O => \N__52313\,
            I => \N__52304\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__52310\,
            I => buf_adcdata_iac_13
        );

    \I__12101\ : Odrv12
    port map (
            O => \N__52307\,
            I => buf_adcdata_iac_13
        );

    \I__12100\ : Odrv4
    port map (
            O => \N__52304\,
            I => buf_adcdata_iac_13
        );

    \I__12099\ : InMux
    port map (
            O => \N__52297\,
            I => \N__52294\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__52294\,
            I => \N__52291\
        );

    \I__12097\ : Span4Mux_h
    port map (
            O => \N__52291\,
            I => \N__52288\
        );

    \I__12096\ : Span4Mux_h
    port map (
            O => \N__52288\,
            I => \N__52285\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__52285\,
            I => n23354
        );

    \I__12094\ : InMux
    port map (
            O => \N__52282\,
            I => \N__52279\
        );

    \I__12093\ : LocalMux
    port map (
            O => \N__52279\,
            I => n23357
        );

    \I__12092\ : InMux
    port map (
            O => \N__52276\,
            I => \N__52273\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__52273\,
            I => \N__52269\
        );

    \I__12090\ : InMux
    port map (
            O => \N__52272\,
            I => \N__52266\
        );

    \I__12089\ : Span4Mux_h
    port map (
            O => \N__52269\,
            I => \N__52263\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__52266\,
            I => data_idxvec_1
        );

    \I__12087\ : Odrv4
    port map (
            O => \N__52263\,
            I => data_idxvec_1
        );

    \I__12086\ : InMux
    port map (
            O => \N__52258\,
            I => \N__52254\
        );

    \I__12085\ : InMux
    port map (
            O => \N__52257\,
            I => \N__52251\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__52254\,
            I => \N__52248\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__52251\,
            I => \N__52242\
        );

    \I__12082\ : Span4Mux_v
    port map (
            O => \N__52248\,
            I => \N__52242\
        );

    \I__12081\ : InMux
    port map (
            O => \N__52247\,
            I => \N__52239\
        );

    \I__12080\ : Odrv4
    port map (
            O => \N__52242\,
            I => data_cntvec_1
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52239\,
            I => data_cntvec_1
        );

    \I__12078\ : InMux
    port map (
            O => \N__52234\,
            I => \N__52230\
        );

    \I__12077\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52226\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__52230\,
            I => \N__52223\
        );

    \I__12075\ : InMux
    port map (
            O => \N__52229\,
            I => \N__52220\
        );

    \I__12074\ : LocalMux
    port map (
            O => \N__52226\,
            I => \N__52215\
        );

    \I__12073\ : Span4Mux_h
    port map (
            O => \N__52223\,
            I => \N__52215\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__52220\,
            I => \N__52212\
        );

    \I__12071\ : Odrv4
    port map (
            O => \N__52215\,
            I => \acadc_skipCount_1\
        );

    \I__12070\ : Odrv4
    port map (
            O => \N__52212\,
            I => \acadc_skipCount_1\
        );

    \I__12069\ : InMux
    port map (
            O => \N__52207\,
            I => \N__52202\
        );

    \I__12068\ : CascadeMux
    port map (
            O => \N__52206\,
            I => \N__52199\
        );

    \I__12067\ : InMux
    port map (
            O => \N__52205\,
            I => \N__52196\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__52202\,
            I => \N__52193\
        );

    \I__12065\ : InMux
    port map (
            O => \N__52199\,
            I => \N__52190\
        );

    \I__12064\ : LocalMux
    port map (
            O => \N__52196\,
            I => req_data_cnt_1
        );

    \I__12063\ : Odrv4
    port map (
            O => \N__52193\,
            I => req_data_cnt_1
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__52190\,
            I => req_data_cnt_1
        );

    \I__12061\ : CascadeMux
    port map (
            O => \N__52183\,
            I => \n22142_cascade_\
        );

    \I__12060\ : InMux
    port map (
            O => \N__52180\,
            I => \N__52177\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__52177\,
            I => \N__52174\
        );

    \I__12058\ : Span4Mux_v
    port map (
            O => \N__52174\,
            I => \N__52171\
        );

    \I__12057\ : Sp12to4
    port map (
            O => \N__52171\,
            I => \N__52168\
        );

    \I__12056\ : Span12Mux_h
    port map (
            O => \N__52168\,
            I => \N__52165\
        );

    \I__12055\ : Odrv12
    port map (
            O => \N__52165\,
            I => n22137
        );

    \I__12054\ : CascadeMux
    port map (
            O => \N__52162\,
            I => \n23408_cascade_\
        );

    \I__12053\ : CascadeMux
    port map (
            O => \N__52159\,
            I => \n23411_cascade_\
        );

    \I__12052\ : InMux
    port map (
            O => \N__52156\,
            I => \N__52153\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__52153\,
            I => \N__52150\
        );

    \I__12050\ : Odrv12
    port map (
            O => \N__52150\,
            I => n111_adj_1754
        );

    \I__12049\ : CascadeMux
    port map (
            O => \N__52147\,
            I => \comm_buf_1_7_N_559_1_cascade_\
        );

    \I__12048\ : InMux
    port map (
            O => \N__52144\,
            I => \N__52139\
        );

    \I__12047\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52135\
        );

    \I__12046\ : CascadeMux
    port map (
            O => \N__52142\,
            I => \N__52131\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__52139\,
            I => \N__52128\
        );

    \I__12044\ : InMux
    port map (
            O => \N__52138\,
            I => \N__52125\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__52135\,
            I => \N__52122\
        );

    \I__12042\ : CascadeMux
    port map (
            O => \N__52134\,
            I => \N__52118\
        );

    \I__12041\ : InMux
    port map (
            O => \N__52131\,
            I => \N__52115\
        );

    \I__12040\ : Span4Mux_v
    port map (
            O => \N__52128\,
            I => \N__52108\
        );

    \I__12039\ : LocalMux
    port map (
            O => \N__52125\,
            I => \N__52108\
        );

    \I__12038\ : Span4Mux_v
    port map (
            O => \N__52122\,
            I => \N__52108\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52121\,
            I => \N__52104\
        );

    \I__12036\ : InMux
    port map (
            O => \N__52118\,
            I => \N__52101\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__52115\,
            I => \N__52098\
        );

    \I__12034\ : Span4Mux_v
    port map (
            O => \N__52108\,
            I => \N__52095\
        );

    \I__12033\ : InMux
    port map (
            O => \N__52107\,
            I => \N__52092\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__52104\,
            I => \N__52087\
        );

    \I__12031\ : LocalMux
    port map (
            O => \N__52101\,
            I => \N__52084\
        );

    \I__12030\ : Span4Mux_v
    port map (
            O => \N__52098\,
            I => \N__52077\
        );

    \I__12029\ : Span4Mux_h
    port map (
            O => \N__52095\,
            I => \N__52077\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__52092\,
            I => \N__52077\
        );

    \I__12027\ : InMux
    port map (
            O => \N__52091\,
            I => \N__52072\
        );

    \I__12026\ : InMux
    port map (
            O => \N__52090\,
            I => \N__52072\
        );

    \I__12025\ : Span4Mux_v
    port map (
            O => \N__52087\,
            I => \N__52069\
        );

    \I__12024\ : Sp12to4
    port map (
            O => \N__52084\,
            I => \N__52066\
        );

    \I__12023\ : Span4Mux_h
    port map (
            O => \N__52077\,
            I => \N__52063\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__52072\,
            I => \N__52060\
        );

    \I__12021\ : Span4Mux_h
    port map (
            O => \N__52069\,
            I => \N__52057\
        );

    \I__12020\ : Span12Mux_v
    port map (
            O => \N__52066\,
            I => \N__52054\
        );

    \I__12019\ : Span4Mux_h
    port map (
            O => \N__52063\,
            I => \N__52051\
        );

    \I__12018\ : Span12Mux_h
    port map (
            O => \N__52060\,
            I => \N__52048\
        );

    \I__12017\ : Odrv4
    port map (
            O => \N__52057\,
            I => comm_buf_1_1
        );

    \I__12016\ : Odrv12
    port map (
            O => \N__52054\,
            I => comm_buf_1_1
        );

    \I__12015\ : Odrv4
    port map (
            O => \N__52051\,
            I => comm_buf_1_1
        );

    \I__12014\ : Odrv12
    port map (
            O => \N__52048\,
            I => comm_buf_1_1
        );

    \I__12013\ : InMux
    port map (
            O => \N__52039\,
            I => \N__52036\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__52036\,
            I => \N__52033\
        );

    \I__12011\ : Span4Mux_h
    port map (
            O => \N__52033\,
            I => \N__52030\
        );

    \I__12010\ : Span4Mux_v
    port map (
            O => \N__52030\,
            I => \N__52027\
        );

    \I__12009\ : Odrv4
    port map (
            O => \N__52027\,
            I => buf_data_iac_9
        );

    \I__12008\ : CascadeMux
    port map (
            O => \N__52024\,
            I => \N__52021\
        );

    \I__12007\ : InMux
    port map (
            O => \N__52021\,
            I => \N__52018\
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__52018\,
            I => n26_adj_1753
        );

    \I__12005\ : InMux
    port map (
            O => \N__52015\,
            I => \N__52012\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__52012\,
            I => n22143
        );

    \I__12003\ : CascadeMux
    port map (
            O => \N__52009\,
            I => \n37_cascade_\
        );

    \I__12002\ : CascadeMux
    port map (
            O => \N__52006\,
            I => \n12761_cascade_\
        );

    \I__12001\ : InMux
    port map (
            O => \N__52003\,
            I => \N__52000\
        );

    \I__12000\ : LocalMux
    port map (
            O => \N__52000\,
            I => \N__51996\
        );

    \I__11999\ : InMux
    port map (
            O => \N__51999\,
            I => \N__51993\
        );

    \I__11998\ : Span4Mux_v
    port map (
            O => \N__51996\,
            I => \N__51990\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__51993\,
            I => data_idxvec_5
        );

    \I__11996\ : Odrv4
    port map (
            O => \N__51990\,
            I => data_idxvec_5
        );

    \I__11995\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51982\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__51982\,
            I => \N__51977\
        );

    \I__11993\ : InMux
    port map (
            O => \N__51981\,
            I => \N__51974\
        );

    \I__11992\ : InMux
    port map (
            O => \N__51980\,
            I => \N__51971\
        );

    \I__11991\ : Span4Mux_h
    port map (
            O => \N__51977\,
            I => \N__51968\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__51974\,
            I => \N__51965\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__51971\,
            I => data_cntvec_5
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__51968\,
            I => data_cntvec_5
        );

    \I__11987\ : Odrv4
    port map (
            O => \N__51965\,
            I => data_cntvec_5
        );

    \I__11986\ : CascadeMux
    port map (
            O => \N__51958\,
            I => \n26_adj_1730_cascade_\
        );

    \I__11985\ : InMux
    port map (
            O => \N__51955\,
            I => \N__51952\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__51952\,
            I => \N__51949\
        );

    \I__11983\ : Span4Mux_v
    port map (
            O => \N__51949\,
            I => \N__51945\
        );

    \I__11982\ : CascadeMux
    port map (
            O => \N__51948\,
            I => \N__51941\
        );

    \I__11981\ : Span4Mux_h
    port map (
            O => \N__51945\,
            I => \N__51938\
        );

    \I__11980\ : InMux
    port map (
            O => \N__51944\,
            I => \N__51933\
        );

    \I__11979\ : InMux
    port map (
            O => \N__51941\,
            I => \N__51933\
        );

    \I__11978\ : Odrv4
    port map (
            O => \N__51938\,
            I => req_data_cnt_5
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__51933\,
            I => req_data_cnt_5
        );

    \I__11976\ : CascadeMux
    port map (
            O => \N__51928\,
            I => \n23336_cascade_\
        );

    \I__11975\ : CascadeMux
    port map (
            O => \N__51925\,
            I => \N__51921\
        );

    \I__11974\ : InMux
    port map (
            O => \N__51924\,
            I => \N__51918\
        );

    \I__11973\ : InMux
    port map (
            O => \N__51921\,
            I => \N__51914\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__51918\,
            I => \N__51911\
        );

    \I__11971\ : InMux
    port map (
            O => \N__51917\,
            I => \N__51908\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__51914\,
            I => \acadc_skipCount_5\
        );

    \I__11969\ : Odrv4
    port map (
            O => \N__51911\,
            I => \acadc_skipCount_5\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__51908\,
            I => \acadc_skipCount_5\
        );

    \I__11967\ : CascadeMux
    port map (
            O => \N__51901\,
            I => \n23339_cascade_\
        );

    \I__11966\ : CascadeMux
    port map (
            O => \N__51898\,
            I => \n30_adj_1731_cascade_\
        );

    \I__11965\ : InMux
    port map (
            O => \N__51895\,
            I => \N__51892\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__51892\,
            I => \N__51889\
        );

    \I__11963\ : Span4Mux_v
    port map (
            O => \N__51889\,
            I => \N__51886\
        );

    \I__11962\ : Span4Mux_h
    port map (
            O => \N__51886\,
            I => \N__51883\
        );

    \I__11961\ : Span4Mux_h
    port map (
            O => \N__51883\,
            I => \N__51880\
        );

    \I__11960\ : Odrv4
    port map (
            O => \N__51880\,
            I => n111_adj_1732
        );

    \I__11959\ : InMux
    port map (
            O => \N__51877\,
            I => \N__51874\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__51874\,
            I => \N__51871\
        );

    \I__11957\ : Span4Mux_h
    port map (
            O => \N__51871\,
            I => \N__51868\
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__51868\,
            I => n22354
        );

    \I__11955\ : CascadeMux
    port map (
            O => \N__51865\,
            I => \N__51862\
        );

    \I__11954\ : InMux
    port map (
            O => \N__51862\,
            I => \N__51859\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__51859\,
            I => n22353
        );

    \I__11952\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51853\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__51853\,
            I => \N__51850\
        );

    \I__11950\ : Span4Mux_h
    port map (
            O => \N__51850\,
            I => \N__51847\
        );

    \I__11949\ : Odrv4
    port map (
            O => \N__51847\,
            I => comm_length_1
        );

    \I__11948\ : InMux
    port map (
            O => \N__51844\,
            I => \N__51841\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__51841\,
            I => n4_adj_1745
        );

    \I__11946\ : InMux
    port map (
            O => \N__51838\,
            I => \N__51834\
        );

    \I__11945\ : InMux
    port map (
            O => \N__51837\,
            I => \N__51831\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__51834\,
            I => \N__51824\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__51831\,
            I => \N__51824\
        );

    \I__11942\ : InMux
    port map (
            O => \N__51830\,
            I => \N__51818\
        );

    \I__11941\ : InMux
    port map (
            O => \N__51829\,
            I => \N__51815\
        );

    \I__11940\ : Span4Mux_v
    port map (
            O => \N__51824\,
            I => \N__51812\
        );

    \I__11939\ : InMux
    port map (
            O => \N__51823\,
            I => \N__51809\
        );

    \I__11938\ : InMux
    port map (
            O => \N__51822\,
            I => \N__51804\
        );

    \I__11937\ : InMux
    port map (
            O => \N__51821\,
            I => \N__51801\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__51818\,
            I => \N__51797\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__51815\,
            I => \N__51792\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__51812\,
            I => \N__51792\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__51809\,
            I => \N__51789\
        );

    \I__11932\ : CascadeMux
    port map (
            O => \N__51808\,
            I => \N__51786\
        );

    \I__11931\ : InMux
    port map (
            O => \N__51807\,
            I => \N__51781\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__51804\,
            I => \N__51774\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51774\
        );

    \I__11928\ : InMux
    port map (
            O => \N__51800\,
            I => \N__51771\
        );

    \I__11927\ : Span4Mux_h
    port map (
            O => \N__51797\,
            I => \N__51768\
        );

    \I__11926\ : Span4Mux_v
    port map (
            O => \N__51792\,
            I => \N__51765\
        );

    \I__11925\ : Span4Mux_h
    port map (
            O => \N__51789\,
            I => \N__51762\
        );

    \I__11924\ : InMux
    port map (
            O => \N__51786\,
            I => \N__51755\
        );

    \I__11923\ : InMux
    port map (
            O => \N__51785\,
            I => \N__51755\
        );

    \I__11922\ : InMux
    port map (
            O => \N__51784\,
            I => \N__51755\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__51781\,
            I => \N__51752\
        );

    \I__11920\ : InMux
    port map (
            O => \N__51780\,
            I => \N__51747\
        );

    \I__11919\ : InMux
    port map (
            O => \N__51779\,
            I => \N__51747\
        );

    \I__11918\ : Odrv12
    port map (
            O => \N__51774\,
            I => comm_index_1
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__51771\,
            I => comm_index_1
        );

    \I__11916\ : Odrv4
    port map (
            O => \N__51768\,
            I => comm_index_1
        );

    \I__11915\ : Odrv4
    port map (
            O => \N__51765\,
            I => comm_index_1
        );

    \I__11914\ : Odrv4
    port map (
            O => \N__51762\,
            I => comm_index_1
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__51755\,
            I => comm_index_1
        );

    \I__11912\ : Odrv4
    port map (
            O => \N__51752\,
            I => comm_index_1
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__51747\,
            I => comm_index_1
        );

    \I__11910\ : InMux
    port map (
            O => \N__51730\,
            I => \N__51726\
        );

    \I__11909\ : CascadeMux
    port map (
            O => \N__51729\,
            I => \N__51722\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__51726\,
            I => \N__51719\
        );

    \I__11907\ : InMux
    port map (
            O => \N__51725\,
            I => \N__51716\
        );

    \I__11906\ : InMux
    port map (
            O => \N__51722\,
            I => \N__51713\
        );

    \I__11905\ : Span4Mux_h
    port map (
            O => \N__51719\,
            I => \N__51708\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__51716\,
            I => \N__51708\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__51713\,
            I => req_data_cnt_14
        );

    \I__11902\ : Odrv4
    port map (
            O => \N__51708\,
            I => req_data_cnt_14
        );

    \I__11901\ : InMux
    port map (
            O => \N__51703\,
            I => \N__51700\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__51700\,
            I => \N__51696\
        );

    \I__11899\ : InMux
    port map (
            O => \N__51699\,
            I => \N__51693\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__51696\,
            I => \N__51690\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__51693\,
            I => data_cntvec_14
        );

    \I__11896\ : Odrv4
    port map (
            O => \N__51690\,
            I => data_cntvec_14
        );

    \I__11895\ : InMux
    port map (
            O => \N__51685\,
            I => \N__51682\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__51682\,
            I => \N__51679\
        );

    \I__11893\ : Span4Mux_h
    port map (
            O => \N__51679\,
            I => \N__51676\
        );

    \I__11892\ : Span4Mux_h
    port map (
            O => \N__51676\,
            I => \N__51673\
        );

    \I__11891\ : Odrv4
    port map (
            O => \N__51673\,
            I => n23
        );

    \I__11890\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51667\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__51667\,
            I => n111
        );

    \I__11888\ : InMux
    port map (
            O => \N__51664\,
            I => \N__51661\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__51661\,
            I => \N__51658\
        );

    \I__11886\ : Odrv4
    port map (
            O => \N__51658\,
            I => n30_adj_1579
        );

    \I__11885\ : InMux
    port map (
            O => \N__51655\,
            I => \N__51652\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__51652\,
            I => \N__51649\
        );

    \I__11883\ : Odrv4
    port map (
            O => \N__51649\,
            I => \comm_buf_1_7_N_559_0\
        );

    \I__11882\ : SRMux
    port map (
            O => \N__51646\,
            I => \N__51642\
        );

    \I__11881\ : SRMux
    port map (
            O => \N__51645\,
            I => \N__51639\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__51642\,
            I => \N__51636\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__51639\,
            I => \N__51633\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__51636\,
            I => \N__51630\
        );

    \I__11877\ : Odrv4
    port map (
            O => \N__51633\,
            I => n21271
        );

    \I__11876\ : Odrv4
    port map (
            O => \N__51630\,
            I => n21271
        );

    \I__11875\ : InMux
    port map (
            O => \N__51625\,
            I => \N__51620\
        );

    \I__11874\ : InMux
    port map (
            O => \N__51624\,
            I => \N__51615\
        );

    \I__11873\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51615\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__51620\,
            I => \N__51609\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__51615\,
            I => \N__51609\
        );

    \I__11870\ : InMux
    port map (
            O => \N__51614\,
            I => \N__51606\
        );

    \I__11869\ : Odrv12
    port map (
            O => \N__51609\,
            I => n11258
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__51606\,
            I => n11258
        );

    \I__11867\ : CascadeMux
    port map (
            O => \N__51601\,
            I => \N__51598\
        );

    \I__11866\ : InMux
    port map (
            O => \N__51598\,
            I => \N__51595\
        );

    \I__11865\ : LocalMux
    port map (
            O => \N__51595\,
            I => \N__51592\
        );

    \I__11864\ : Odrv4
    port map (
            O => \N__51592\,
            I => n22089
        );

    \I__11863\ : InMux
    port map (
            O => \N__51589\,
            I => \N__51586\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__51586\,
            I => \N__51582\
        );

    \I__11861\ : InMux
    port map (
            O => \N__51585\,
            I => \N__51579\
        );

    \I__11860\ : Odrv4
    port map (
            O => \N__51582\,
            I => n20318
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__51579\,
            I => n20318
        );

    \I__11858\ : CascadeMux
    port map (
            O => \N__51574\,
            I => \n12_adj_1677_cascade_\
        );

    \I__11857\ : CascadeMux
    port map (
            O => \N__51571\,
            I => \n12892_cascade_\
        );

    \I__11856\ : InMux
    port map (
            O => \N__51568\,
            I => \N__51563\
        );

    \I__11855\ : InMux
    port map (
            O => \N__51567\,
            I => \N__51560\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51566\,
            I => \N__51557\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__51563\,
            I => \N__51554\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__51560\,
            I => n12951
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__51557\,
            I => n12951
        );

    \I__11850\ : Odrv4
    port map (
            O => \N__51554\,
            I => n12951
        );

    \I__11849\ : CascadeMux
    port map (
            O => \N__51547\,
            I => \N__51543\
        );

    \I__11848\ : CascadeMux
    port map (
            O => \N__51546\,
            I => \N__51539\
        );

    \I__11847\ : InMux
    port map (
            O => \N__51543\,
            I => \N__51536\
        );

    \I__11846\ : InMux
    port map (
            O => \N__51542\,
            I => \N__51531\
        );

    \I__11845\ : InMux
    port map (
            O => \N__51539\,
            I => \N__51531\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__51536\,
            I => \N__51528\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__51531\,
            I => \N__51525\
        );

    \I__11842\ : Span12Mux_v
    port map (
            O => \N__51528\,
            I => \N__51522\
        );

    \I__11841\ : Span12Mux_v
    port map (
            O => \N__51525\,
            I => \N__51519\
        );

    \I__11840\ : Odrv12
    port map (
            O => \N__51522\,
            I => n9714
        );

    \I__11839\ : Odrv12
    port map (
            O => \N__51519\,
            I => n9714
        );

    \I__11838\ : InMux
    port map (
            O => \N__51514\,
            I => \N__51511\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__51511\,
            I => \N__51508\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__51508\,
            I => \N__51505\
        );

    \I__11835\ : Odrv4
    port map (
            O => \N__51505\,
            I => n11_adj_1585
        );

    \I__11834\ : InMux
    port map (
            O => \N__51502\,
            I => \N__51498\
        );

    \I__11833\ : InMux
    port map (
            O => \N__51501\,
            I => \N__51495\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__51498\,
            I => \N__51492\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__51495\,
            I => \N__51489\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__51492\,
            I => \N__51486\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__51489\,
            I => \N__51483\
        );

    \I__11828\ : Span4Mux_h
    port map (
            O => \N__51486\,
            I => \N__51478\
        );

    \I__11827\ : Span4Mux_v
    port map (
            O => \N__51483\,
            I => \N__51478\
        );

    \I__11826\ : Span4Mux_v
    port map (
            O => \N__51478\,
            I => \N__51475\
        );

    \I__11825\ : Odrv4
    port map (
            O => \N__51475\,
            I => n14_adj_1652
        );

    \I__11824\ : InMux
    port map (
            O => \N__51472\,
            I => \N__51462\
        );

    \I__11823\ : InMux
    port map (
            O => \N__51471\,
            I => \N__51462\
        );

    \I__11822\ : InMux
    port map (
            O => \N__51470\,
            I => \N__51462\
        );

    \I__11821\ : InMux
    port map (
            O => \N__51469\,
            I => \N__51459\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__51462\,
            I => \N__51454\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__51459\,
            I => \N__51454\
        );

    \I__11818\ : Odrv4
    port map (
            O => \N__51454\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__11817\ : CascadeMux
    port map (
            O => \N__51451\,
            I => \N__51447\
        );

    \I__11816\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51441\
        );

    \I__11815\ : InMux
    port map (
            O => \N__51447\,
            I => \N__51432\
        );

    \I__11814\ : InMux
    port map (
            O => \N__51446\,
            I => \N__51432\
        );

    \I__11813\ : InMux
    port map (
            O => \N__51445\,
            I => \N__51432\
        );

    \I__11812\ : InMux
    port map (
            O => \N__51444\,
            I => \N__51432\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__51441\,
            I => \N__51429\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__51432\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__11809\ : Odrv4
    port map (
            O => \N__51429\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__11808\ : InMux
    port map (
            O => \N__51424\,
            I => \N__51417\
        );

    \I__11807\ : InMux
    port map (
            O => \N__51423\,
            I => \N__51417\
        );

    \I__11806\ : InMux
    port map (
            O => \N__51422\,
            I => \N__51414\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__51417\,
            I => \N__51409\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__51414\,
            I => \N__51409\
        );

    \I__11803\ : Odrv4
    port map (
            O => \N__51409\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__11802\ : InMux
    port map (
            O => \N__51406\,
            I => \N__51403\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__51403\,
            I => \N__51400\
        );

    \I__11800\ : Odrv4
    port map (
            O => \N__51400\,
            I => n22487
        );

    \I__11799\ : InMux
    port map (
            O => \N__51397\,
            I => \N__51393\
        );

    \I__11798\ : InMux
    port map (
            O => \N__51396\,
            I => \N__51390\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__51393\,
            I => \N__51387\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__51390\,
            I => \N__51384\
        );

    \I__11795\ : Span4Mux_h
    port map (
            O => \N__51387\,
            I => \N__51381\
        );

    \I__11794\ : Span12Mux_h
    port map (
            O => \N__51384\,
            I => \N__51377\
        );

    \I__11793\ : Span4Mux_h
    port map (
            O => \N__51381\,
            I => \N__51374\
        );

    \I__11792\ : InMux
    port map (
            O => \N__51380\,
            I => \N__51371\
        );

    \I__11791\ : Odrv12
    port map (
            O => \N__51377\,
            I => n21983
        );

    \I__11790\ : Odrv4
    port map (
            O => \N__51374\,
            I => n21983
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__51371\,
            I => n21983
        );

    \I__11788\ : InMux
    port map (
            O => \N__51364\,
            I => \N__51355\
        );

    \I__11787\ : InMux
    port map (
            O => \N__51363\,
            I => \N__51355\
        );

    \I__11786\ : InMux
    port map (
            O => \N__51362\,
            I => \N__51349\
        );

    \I__11785\ : InMux
    port map (
            O => \N__51361\,
            I => \N__51343\
        );

    \I__11784\ : InMux
    port map (
            O => \N__51360\,
            I => \N__51343\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__51355\,
            I => \N__51340\
        );

    \I__11782\ : InMux
    port map (
            O => \N__51354\,
            I => \N__51331\
        );

    \I__11781\ : InMux
    port map (
            O => \N__51353\,
            I => \N__51331\
        );

    \I__11780\ : InMux
    port map (
            O => \N__51352\,
            I => \N__51331\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__51349\,
            I => \N__51328\
        );

    \I__11778\ : InMux
    port map (
            O => \N__51348\,
            I => \N__51325\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__51343\,
            I => \N__51320\
        );

    \I__11776\ : Span4Mux_v
    port map (
            O => \N__51340\,
            I => \N__51317\
        );

    \I__11775\ : InMux
    port map (
            O => \N__51339\,
            I => \N__51314\
        );

    \I__11774\ : CascadeMux
    port map (
            O => \N__51338\,
            I => \N__51311\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51331\,
            I => \N__51307\
        );

    \I__11772\ : Span4Mux_h
    port map (
            O => \N__51328\,
            I => \N__51302\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__51325\,
            I => \N__51302\
        );

    \I__11770\ : InMux
    port map (
            O => \N__51324\,
            I => \N__51299\
        );

    \I__11769\ : InMux
    port map (
            O => \N__51323\,
            I => \N__51296\
        );

    \I__11768\ : Span4Mux_v
    port map (
            O => \N__51320\,
            I => \N__51289\
        );

    \I__11767\ : Span4Mux_h
    port map (
            O => \N__51317\,
            I => \N__51289\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__51314\,
            I => \N__51289\
        );

    \I__11765\ : InMux
    port map (
            O => \N__51311\,
            I => \N__51284\
        );

    \I__11764\ : InMux
    port map (
            O => \N__51310\,
            I => \N__51284\
        );

    \I__11763\ : Span4Mux_v
    port map (
            O => \N__51307\,
            I => \N__51280\
        );

    \I__11762\ : Span4Mux_h
    port map (
            O => \N__51302\,
            I => \N__51277\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__51299\,
            I => \N__51268\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__51296\,
            I => \N__51268\
        );

    \I__11759\ : Span4Mux_h
    port map (
            O => \N__51289\,
            I => \N__51268\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__51284\,
            I => \N__51268\
        );

    \I__11757\ : InMux
    port map (
            O => \N__51283\,
            I => \N__51265\
        );

    \I__11756\ : Span4Mux_h
    port map (
            O => \N__51280\,
            I => \N__51262\
        );

    \I__11755\ : Span4Mux_h
    port map (
            O => \N__51277\,
            I => \N__51259\
        );

    \I__11754\ : Span4Mux_v
    port map (
            O => \N__51268\,
            I => \N__51256\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__51265\,
            I => n13171
        );

    \I__11752\ : Odrv4
    port map (
            O => \N__51262\,
            I => n13171
        );

    \I__11751\ : Odrv4
    port map (
            O => \N__51259\,
            I => n13171
        );

    \I__11750\ : Odrv4
    port map (
            O => \N__51256\,
            I => n13171
        );

    \I__11749\ : CascadeMux
    port map (
            O => \N__51247\,
            I => \n13171_cascade_\
        );

    \I__11748\ : InMux
    port map (
            O => \N__51244\,
            I => \N__51241\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51241\,
            I => n22033
        );

    \I__11746\ : CascadeMux
    port map (
            O => \N__51238\,
            I => \n12064_cascade_\
        );

    \I__11745\ : CEMux
    port map (
            O => \N__51235\,
            I => \N__51232\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__51232\,
            I => n21885
        );

    \I__11743\ : CascadeMux
    port map (
            O => \N__51229\,
            I => \n22073_cascade_\
        );

    \I__11742\ : SRMux
    port map (
            O => \N__51226\,
            I => \N__51220\
        );

    \I__11741\ : SRMux
    port map (
            O => \N__51225\,
            I => \N__51216\
        );

    \I__11740\ : SRMux
    port map (
            O => \N__51224\,
            I => \N__51213\
        );

    \I__11739\ : SRMux
    port map (
            O => \N__51223\,
            I => \N__51210\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__51220\,
            I => \N__51207\
        );

    \I__11737\ : SRMux
    port map (
            O => \N__51219\,
            I => \N__51204\
        );

    \I__11736\ : LocalMux
    port map (
            O => \N__51216\,
            I => \N__51197\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__51213\,
            I => \N__51197\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__51210\,
            I => \N__51197\
        );

    \I__11733\ : Span4Mux_v
    port map (
            O => \N__51207\,
            I => \N__51192\
        );

    \I__11732\ : LocalMux
    port map (
            O => \N__51204\,
            I => \N__51192\
        );

    \I__11731\ : Span4Mux_v
    port map (
            O => \N__51197\,
            I => \N__51189\
        );

    \I__11730\ : Odrv4
    port map (
            O => \N__51192\,
            I => flagcntwd
        );

    \I__11729\ : Odrv4
    port map (
            O => \N__51189\,
            I => flagcntwd
        );

    \I__11728\ : CEMux
    port map (
            O => \N__51184\,
            I => \N__51181\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__51181\,
            I => \N__51178\
        );

    \I__11726\ : Odrv4
    port map (
            O => \N__51178\,
            I => n12050
        );

    \I__11725\ : InMux
    port map (
            O => \N__51175\,
            I => \N__51172\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__51172\,
            I => n10_adj_1602
        );

    \I__11723\ : InMux
    port map (
            O => \N__51169\,
            I => \N__51161\
        );

    \I__11722\ : InMux
    port map (
            O => \N__51168\,
            I => \N__51158\
        );

    \I__11721\ : InMux
    port map (
            O => \N__51167\,
            I => \N__51153\
        );

    \I__11720\ : InMux
    port map (
            O => \N__51166\,
            I => \N__51153\
        );

    \I__11719\ : InMux
    port map (
            O => \N__51165\,
            I => \N__51148\
        );

    \I__11718\ : InMux
    port map (
            O => \N__51164\,
            I => \N__51148\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__51161\,
            I => \N__51141\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__51158\,
            I => \N__51141\
        );

    \I__11715\ : LocalMux
    port map (
            O => \N__51153\,
            I => \N__51141\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__51148\,
            I => \N__51136\
        );

    \I__11713\ : Span4Mux_v
    port map (
            O => \N__51141\,
            I => \N__51136\
        );

    \I__11712\ : Odrv4
    port map (
            O => \N__51136\,
            I => comm_cmd_7
        );

    \I__11711\ : CascadeMux
    port map (
            O => \N__51133\,
            I => \N__51130\
        );

    \I__11710\ : InMux
    port map (
            O => \N__51130\,
            I => \N__51127\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__51127\,
            I => n29
        );

    \I__11708\ : InMux
    port map (
            O => \N__51124\,
            I => \N__51121\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__51121\,
            I => \N__51118\
        );

    \I__11706\ : Span4Mux_v
    port map (
            O => \N__51118\,
            I => \N__51115\
        );

    \I__11705\ : Span4Mux_h
    port map (
            O => \N__51115\,
            I => \N__51111\
        );

    \I__11704\ : InMux
    port map (
            O => \N__51114\,
            I => \N__51108\
        );

    \I__11703\ : Odrv4
    port map (
            O => \N__51111\,
            I => \comm_spi.n24034\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__51108\,
            I => \comm_spi.n24034\
        );

    \I__11701\ : InMux
    port map (
            O => \N__51103\,
            I => \N__51100\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__51100\,
            I => \N__51097\
        );

    \I__11699\ : Span4Mux_h
    port map (
            O => \N__51097\,
            I => \N__51094\
        );

    \I__11698\ : Span4Mux_h
    port map (
            O => \N__51094\,
            I => \N__51090\
        );

    \I__11697\ : InMux
    port map (
            O => \N__51093\,
            I => \N__51087\
        );

    \I__11696\ : Sp12to4
    port map (
            O => \N__51090\,
            I => \N__51082\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__51087\,
            I => \N__51082\
        );

    \I__11694\ : Odrv12
    port map (
            O => \N__51082\,
            I => \comm_spi.n15352\
        );

    \I__11693\ : InMux
    port map (
            O => \N__51079\,
            I => \N__51076\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__51076\,
            I => \N__51072\
        );

    \I__11691\ : InMux
    port map (
            O => \N__51075\,
            I => \N__51069\
        );

    \I__11690\ : Span4Mux_h
    port map (
            O => \N__51072\,
            I => \N__51066\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__51069\,
            I => \N__51063\
        );

    \I__11688\ : Span4Mux_h
    port map (
            O => \N__51066\,
            I => \N__51060\
        );

    \I__11687\ : Span4Mux_v
    port map (
            O => \N__51063\,
            I => \N__51057\
        );

    \I__11686\ : Odrv4
    port map (
            O => \N__51060\,
            I => \comm_spi.n15353\
        );

    \I__11685\ : Odrv4
    port map (
            O => \N__51057\,
            I => \comm_spi.n15353\
        );

    \I__11684\ : InMux
    port map (
            O => \N__51052\,
            I => \N__51049\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__51049\,
            I => \N__51046\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__51046\,
            I => \N__51042\
        );

    \I__11681\ : InMux
    port map (
            O => \N__51045\,
            I => \N__51039\
        );

    \I__11680\ : Span4Mux_v
    port map (
            O => \N__51042\,
            I => \N__51036\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__51039\,
            I => \N__51033\
        );

    \I__11678\ : Span4Mux_h
    port map (
            O => \N__51036\,
            I => \N__51028\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__51033\,
            I => \N__51028\
        );

    \I__11676\ : Span4Mux_h
    port map (
            O => \N__51028\,
            I => \N__51025\
        );

    \I__11675\ : Odrv4
    port map (
            O => \N__51025\,
            I => \comm_spi.n15357\
        );

    \I__11674\ : SRMux
    port map (
            O => \N__51022\,
            I => \N__51019\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__51019\,
            I => \N__51016\
        );

    \I__11672\ : Span4Mux_v
    port map (
            O => \N__51016\,
            I => \N__51013\
        );

    \I__11671\ : Span4Mux_h
    port map (
            O => \N__51013\,
            I => \N__51010\
        );

    \I__11670\ : Span4Mux_v
    port map (
            O => \N__51010\,
            I => \N__51007\
        );

    \I__11669\ : Odrv4
    port map (
            O => \N__51007\,
            I => \comm_spi.data_tx_7__N_874\
        );

    \I__11668\ : CascadeMux
    port map (
            O => \N__51004\,
            I => \n22489_cascade_\
        );

    \I__11667\ : CascadeMux
    port map (
            O => \N__51001\,
            I => \n20959_cascade_\
        );

    \I__11666\ : CEMux
    port map (
            O => \N__50998\,
            I => \N__50995\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__50995\,
            I => n21883
        );

    \I__11664\ : InMux
    port map (
            O => \N__50992\,
            I => \N__50989\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__50989\,
            I => n19241
        );

    \I__11662\ : InMux
    port map (
            O => \N__50986\,
            I => \N__50983\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__50983\,
            I => \N__50980\
        );

    \I__11660\ : Odrv12
    port map (
            O => \N__50980\,
            I => n22177
        );

    \I__11659\ : InMux
    port map (
            O => \N__50977\,
            I => \N__50974\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__50974\,
            I => \N__50971\
        );

    \I__11657\ : Odrv12
    port map (
            O => \N__50971\,
            I => n22180
        );

    \I__11656\ : CascadeMux
    port map (
            O => \N__50968\,
            I => \n23462_cascade_\
        );

    \I__11655\ : InMux
    port map (
            O => \N__50965\,
            I => \N__50962\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__50962\,
            I => \N__50959\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__50959\,
            I => \N__50956\
        );

    \I__11652\ : Odrv4
    port map (
            O => \N__50956\,
            I => n23465
        );

    \I__11651\ : CascadeMux
    port map (
            O => \N__50953\,
            I => \N__50950\
        );

    \I__11650\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50946\
        );

    \I__11649\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50943\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__50946\,
            I => data_idxvec_9
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__50943\,
            I => data_idxvec_9
        );

    \I__11646\ : InMux
    port map (
            O => \N__50938\,
            I => \N__50934\
        );

    \I__11645\ : InMux
    port map (
            O => \N__50937\,
            I => \N__50930\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__50934\,
            I => \N__50927\
        );

    \I__11643\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50924\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__50930\,
            I => data_cntvec_9
        );

    \I__11641\ : Odrv4
    port map (
            O => \N__50927\,
            I => data_cntvec_9
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__50924\,
            I => data_cntvec_9
        );

    \I__11639\ : InMux
    port map (
            O => \N__50917\,
            I => \N__50914\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__50914\,
            I => \N__50911\
        );

    \I__11637\ : Span4Mux_v
    port map (
            O => \N__50911\,
            I => \N__50908\
        );

    \I__11636\ : Span4Mux_h
    port map (
            O => \N__50908\,
            I => \N__50905\
        );

    \I__11635\ : Odrv4
    port map (
            O => \N__50905\,
            I => buf_data_iac_17
        );

    \I__11634\ : CascadeMux
    port map (
            O => \N__50902\,
            I => \n22184_cascade_\
        );

    \I__11633\ : InMux
    port map (
            O => \N__50899\,
            I => \N__50896\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__50896\,
            I => n22186
        );

    \I__11631\ : InMux
    port map (
            O => \N__50893\,
            I => \N__50880\
        );

    \I__11630\ : InMux
    port map (
            O => \N__50892\,
            I => \N__50880\
        );

    \I__11629\ : InMux
    port map (
            O => \N__50891\,
            I => \N__50877\
        );

    \I__11628\ : InMux
    port map (
            O => \N__50890\,
            I => \N__50872\
        );

    \I__11627\ : InMux
    port map (
            O => \N__50889\,
            I => \N__50872\
        );

    \I__11626\ : InMux
    port map (
            O => \N__50888\,
            I => \N__50865\
        );

    \I__11625\ : InMux
    port map (
            O => \N__50887\,
            I => \N__50865\
        );

    \I__11624\ : InMux
    port map (
            O => \N__50886\,
            I => \N__50865\
        );

    \I__11623\ : CascadeMux
    port map (
            O => \N__50885\,
            I => \N__50862\
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__50880\,
            I => \N__50859\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__50877\,
            I => \N__50853\
        );

    \I__11620\ : LocalMux
    port map (
            O => \N__50872\,
            I => \N__50853\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__50865\,
            I => \N__50850\
        );

    \I__11618\ : InMux
    port map (
            O => \N__50862\,
            I => \N__50847\
        );

    \I__11617\ : Span4Mux_h
    port map (
            O => \N__50859\,
            I => \N__50844\
        );

    \I__11616\ : InMux
    port map (
            O => \N__50858\,
            I => \N__50841\
        );

    \I__11615\ : Span4Mux_v
    port map (
            O => \N__50853\,
            I => \N__50836\
        );

    \I__11614\ : Span4Mux_h
    port map (
            O => \N__50850\,
            I => \N__50836\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__50847\,
            I => \N__50833\
        );

    \I__11612\ : Span4Mux_h
    port map (
            O => \N__50844\,
            I => \N__50828\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__50841\,
            I => \N__50828\
        );

    \I__11610\ : Span4Mux_h
    port map (
            O => \N__50836\,
            I => \N__50825\
        );

    \I__11609\ : Span12Mux_s11_h
    port map (
            O => \N__50833\,
            I => \N__50820\
        );

    \I__11608\ : Sp12to4
    port map (
            O => \N__50828\,
            I => \N__50820\
        );

    \I__11607\ : Odrv4
    port map (
            O => \N__50825\,
            I => n21997
        );

    \I__11606\ : Odrv12
    port map (
            O => \N__50820\,
            I => n21997
        );

    \I__11605\ : InMux
    port map (
            O => \N__50815\,
            I => \N__50809\
        );

    \I__11604\ : InMux
    port map (
            O => \N__50814\,
            I => \N__50809\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__50809\,
            I => \N__50804\
        );

    \I__11602\ : InMux
    port map (
            O => \N__50808\,
            I => \N__50801\
        );

    \I__11601\ : InMux
    port map (
            O => \N__50807\,
            I => \N__50798\
        );

    \I__11600\ : Span4Mux_v
    port map (
            O => \N__50804\,
            I => \N__50794\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__50801\,
            I => \N__50791\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__50798\,
            I => \N__50788\
        );

    \I__11597\ : InMux
    port map (
            O => \N__50797\,
            I => \N__50785\
        );

    \I__11596\ : Odrv4
    port map (
            O => \N__50794\,
            I => n14_adj_1656
        );

    \I__11595\ : Odrv12
    port map (
            O => \N__50791\,
            I => n14_adj_1656
        );

    \I__11594\ : Odrv4
    port map (
            O => \N__50788\,
            I => n14_adj_1656
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__50785\,
            I => n14_adj_1656
        );

    \I__11592\ : InMux
    port map (
            O => \N__50776\,
            I => \N__50772\
        );

    \I__11591\ : InMux
    port map (
            O => \N__50775\,
            I => \N__50765\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__50772\,
            I => \N__50760\
        );

    \I__11589\ : InMux
    port map (
            O => \N__50771\,
            I => \N__50755\
        );

    \I__11588\ : InMux
    port map (
            O => \N__50770\,
            I => \N__50755\
        );

    \I__11587\ : InMux
    port map (
            O => \N__50769\,
            I => \N__50748\
        );

    \I__11586\ : InMux
    port map (
            O => \N__50768\,
            I => \N__50748\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__50765\,
            I => \N__50745\
        );

    \I__11584\ : InMux
    port map (
            O => \N__50764\,
            I => \N__50742\
        );

    \I__11583\ : InMux
    port map (
            O => \N__50763\,
            I => \N__50739\
        );

    \I__11582\ : Span4Mux_v
    port map (
            O => \N__50760\,
            I => \N__50733\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__50755\,
            I => \N__50730\
        );

    \I__11580\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50727\
        );

    \I__11579\ : InMux
    port map (
            O => \N__50753\,
            I => \N__50724\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__50748\,
            I => \N__50719\
        );

    \I__11577\ : Span4Mux_v
    port map (
            O => \N__50745\,
            I => \N__50716\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__50742\,
            I => \N__50711\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__50739\,
            I => \N__50711\
        );

    \I__11574\ : InMux
    port map (
            O => \N__50738\,
            I => \N__50704\
        );

    \I__11573\ : InMux
    port map (
            O => \N__50737\,
            I => \N__50704\
        );

    \I__11572\ : InMux
    port map (
            O => \N__50736\,
            I => \N__50704\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__50733\,
            I => \N__50697\
        );

    \I__11570\ : Span4Mux_v
    port map (
            O => \N__50730\,
            I => \N__50697\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__50727\,
            I => \N__50697\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__50724\,
            I => \N__50694\
        );

    \I__11567\ : InMux
    port map (
            O => \N__50723\,
            I => \N__50689\
        );

    \I__11566\ : InMux
    port map (
            O => \N__50722\,
            I => \N__50689\
        );

    \I__11565\ : Span4Mux_v
    port map (
            O => \N__50719\,
            I => \N__50685\
        );

    \I__11564\ : Span4Mux_h
    port map (
            O => \N__50716\,
            I => \N__50682\
        );

    \I__11563\ : Span4Mux_v
    port map (
            O => \N__50711\,
            I => \N__50679\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__50704\,
            I => \N__50676\
        );

    \I__11561\ : Span4Mux_v
    port map (
            O => \N__50697\,
            I => \N__50669\
        );

    \I__11560\ : Span4Mux_h
    port map (
            O => \N__50694\,
            I => \N__50669\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__50689\,
            I => \N__50669\
        );

    \I__11558\ : InMux
    port map (
            O => \N__50688\,
            I => \N__50666\
        );

    \I__11557\ : Span4Mux_h
    port map (
            O => \N__50685\,
            I => \N__50659\
        );

    \I__11556\ : Span4Mux_v
    port map (
            O => \N__50682\,
            I => \N__50659\
        );

    \I__11555\ : Span4Mux_h
    port map (
            O => \N__50679\,
            I => \N__50659\
        );

    \I__11554\ : Span12Mux_v
    port map (
            O => \N__50676\,
            I => \N__50656\
        );

    \I__11553\ : Span4Mux_v
    port map (
            O => \N__50669\,
            I => \N__50653\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__50666\,
            I => n13093
        );

    \I__11551\ : Odrv4
    port map (
            O => \N__50659\,
            I => n13093
        );

    \I__11550\ : Odrv12
    port map (
            O => \N__50656\,
            I => n13093
        );

    \I__11549\ : Odrv4
    port map (
            O => \N__50653\,
            I => n13093
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__50644\,
            I => \N__50641\
        );

    \I__11547\ : InMux
    port map (
            O => \N__50641\,
            I => \N__50637\
        );

    \I__11546\ : InMux
    port map (
            O => \N__50640\,
            I => \N__50634\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__50637\,
            I => \N__50630\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__50634\,
            I => \N__50627\
        );

    \I__11543\ : InMux
    port map (
            O => \N__50633\,
            I => \N__50624\
        );

    \I__11542\ : Span12Mux_h
    port map (
            O => \N__50630\,
            I => \N__50621\
        );

    \I__11541\ : Odrv12
    port map (
            O => \N__50627\,
            I => buf_dds0_9
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__50624\,
            I => buf_dds0_9
        );

    \I__11539\ : Odrv12
    port map (
            O => \N__50621\,
            I => buf_dds0_9
        );

    \I__11538\ : InMux
    port map (
            O => \N__50614\,
            I => \N__50611\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__50611\,
            I => \N__50605\
        );

    \I__11536\ : InMux
    port map (
            O => \N__50610\,
            I => \N__50600\
        );

    \I__11535\ : InMux
    port map (
            O => \N__50609\,
            I => \N__50600\
        );

    \I__11534\ : InMux
    port map (
            O => \N__50608\,
            I => \N__50596\
        );

    \I__11533\ : Span4Mux_h
    port map (
            O => \N__50605\,
            I => \N__50587\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__50600\,
            I => \N__50587\
        );

    \I__11531\ : InMux
    port map (
            O => \N__50599\,
            I => \N__50584\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__50596\,
            I => \N__50581\
        );

    \I__11529\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50578\
        );

    \I__11528\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50573\
        );

    \I__11527\ : InMux
    port map (
            O => \N__50593\,
            I => \N__50573\
        );

    \I__11526\ : InMux
    port map (
            O => \N__50592\,
            I => \N__50570\
        );

    \I__11525\ : Span4Mux_h
    port map (
            O => \N__50587\,
            I => \N__50567\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__50584\,
            I => dds_state_0
        );

    \I__11523\ : Odrv4
    port map (
            O => \N__50581\,
            I => dds_state_0
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__50578\,
            I => dds_state_0
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__50573\,
            I => dds_state_0
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__50570\,
            I => dds_state_0
        );

    \I__11519\ : Odrv4
    port map (
            O => \N__50567\,
            I => dds_state_0
        );

    \I__11518\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50532\
        );

    \I__11517\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50521\
        );

    \I__11516\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50521\
        );

    \I__11515\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50521\
        );

    \I__11514\ : InMux
    port map (
            O => \N__50550\,
            I => \N__50521\
        );

    \I__11513\ : InMux
    port map (
            O => \N__50549\,
            I => \N__50521\
        );

    \I__11512\ : InMux
    port map (
            O => \N__50548\,
            I => \N__50510\
        );

    \I__11511\ : InMux
    port map (
            O => \N__50547\,
            I => \N__50510\
        );

    \I__11510\ : InMux
    port map (
            O => \N__50546\,
            I => \N__50510\
        );

    \I__11509\ : InMux
    port map (
            O => \N__50545\,
            I => \N__50510\
        );

    \I__11508\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50510\
        );

    \I__11507\ : InMux
    port map (
            O => \N__50543\,
            I => \N__50507\
        );

    \I__11506\ : InMux
    port map (
            O => \N__50542\,
            I => \N__50498\
        );

    \I__11505\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50498\
        );

    \I__11504\ : InMux
    port map (
            O => \N__50540\,
            I => \N__50498\
        );

    \I__11503\ : InMux
    port map (
            O => \N__50539\,
            I => \N__50498\
        );

    \I__11502\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50495\
        );

    \I__11501\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50492\
        );

    \I__11500\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50485\
        );

    \I__11499\ : InMux
    port map (
            O => \N__50535\,
            I => \N__50485\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__50532\,
            I => \N__50480\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__50521\,
            I => \N__50480\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__50510\,
            I => \N__50477\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__50507\,
            I => \N__50474\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__50498\,
            I => \N__50471\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__50495\,
            I => \N__50466\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__50492\,
            I => \N__50466\
        );

    \I__11491\ : InMux
    port map (
            O => \N__50491\,
            I => \N__50461\
        );

    \I__11490\ : InMux
    port map (
            O => \N__50490\,
            I => \N__50461\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__50485\,
            I => \N__50456\
        );

    \I__11488\ : Span4Mux_h
    port map (
            O => \N__50480\,
            I => \N__50452\
        );

    \I__11487\ : Span12Mux_v
    port map (
            O => \N__50477\,
            I => \N__50449\
        );

    \I__11486\ : Span4Mux_h
    port map (
            O => \N__50474\,
            I => \N__50440\
        );

    \I__11485\ : Span4Mux_v
    port map (
            O => \N__50471\,
            I => \N__50440\
        );

    \I__11484\ : Span4Mux_v
    port map (
            O => \N__50466\,
            I => \N__50440\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__50461\,
            I => \N__50440\
        );

    \I__11482\ : InMux
    port map (
            O => \N__50460\,
            I => \N__50435\
        );

    \I__11481\ : InMux
    port map (
            O => \N__50459\,
            I => \N__50435\
        );

    \I__11480\ : Span4Mux_h
    port map (
            O => \N__50456\,
            I => \N__50432\
        );

    \I__11479\ : InMux
    port map (
            O => \N__50455\,
            I => \N__50429\
        );

    \I__11478\ : Odrv4
    port map (
            O => \N__50452\,
            I => dds_state_2
        );

    \I__11477\ : Odrv12
    port map (
            O => \N__50449\,
            I => dds_state_2
        );

    \I__11476\ : Odrv4
    port map (
            O => \N__50440\,
            I => dds_state_2
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__50435\,
            I => dds_state_2
        );

    \I__11474\ : Odrv4
    port map (
            O => \N__50432\,
            I => dds_state_2
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__50429\,
            I => dds_state_2
        );

    \I__11472\ : InMux
    port map (
            O => \N__50416\,
            I => \N__50390\
        );

    \I__11471\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50390\
        );

    \I__11470\ : InMux
    port map (
            O => \N__50414\,
            I => \N__50390\
        );

    \I__11469\ : InMux
    port map (
            O => \N__50413\,
            I => \N__50390\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50412\,
            I => \N__50390\
        );

    \I__11467\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50390\
        );

    \I__11466\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50379\
        );

    \I__11465\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50379\
        );

    \I__11464\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50379\
        );

    \I__11463\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50379\
        );

    \I__11462\ : InMux
    port map (
            O => \N__50406\,
            I => \N__50379\
        );

    \I__11461\ : SRMux
    port map (
            O => \N__50405\,
            I => \N__50376\
        );

    \I__11460\ : CEMux
    port map (
            O => \N__50404\,
            I => \N__50369\
        );

    \I__11459\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50365\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__50390\,
            I => \N__50360\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__50379\,
            I => \N__50357\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__50376\,
            I => \N__50354\
        );

    \I__11455\ : InMux
    port map (
            O => \N__50375\,
            I => \N__50345\
        );

    \I__11454\ : InMux
    port map (
            O => \N__50374\,
            I => \N__50345\
        );

    \I__11453\ : InMux
    port map (
            O => \N__50373\,
            I => \N__50345\
        );

    \I__11452\ : InMux
    port map (
            O => \N__50372\,
            I => \N__50345\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__50369\,
            I => \N__50342\
        );

    \I__11450\ : InMux
    port map (
            O => \N__50368\,
            I => \N__50339\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__50365\,
            I => \N__50336\
        );

    \I__11448\ : InMux
    port map (
            O => \N__50364\,
            I => \N__50331\
        );

    \I__11447\ : InMux
    port map (
            O => \N__50363\,
            I => \N__50331\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__50360\,
            I => \N__50326\
        );

    \I__11445\ : Span4Mux_h
    port map (
            O => \N__50357\,
            I => \N__50319\
        );

    \I__11444\ : Span4Mux_h
    port map (
            O => \N__50354\,
            I => \N__50319\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__50345\,
            I => \N__50319\
        );

    \I__11442\ : Span4Mux_v
    port map (
            O => \N__50342\,
            I => \N__50311\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__50339\,
            I => \N__50304\
        );

    \I__11440\ : Span4Mux_h
    port map (
            O => \N__50336\,
            I => \N__50304\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__50331\,
            I => \N__50304\
        );

    \I__11438\ : InMux
    port map (
            O => \N__50330\,
            I => \N__50301\
        );

    \I__11437\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50298\
        );

    \I__11436\ : Span4Mux_h
    port map (
            O => \N__50326\,
            I => \N__50293\
        );

    \I__11435\ : Span4Mux_h
    port map (
            O => \N__50319\,
            I => \N__50293\
        );

    \I__11434\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50288\
        );

    \I__11433\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50288\
        );

    \I__11432\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50281\
        );

    \I__11431\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50281\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50314\,
            I => \N__50281\
        );

    \I__11429\ : Span4Mux_h
    port map (
            O => \N__50311\,
            I => \N__50276\
        );

    \I__11428\ : Span4Mux_h
    port map (
            O => \N__50304\,
            I => \N__50276\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__50301\,
            I => dds_state_1
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__50298\,
            I => dds_state_1
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__50293\,
            I => dds_state_1
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__50288\,
            I => dds_state_1
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__50281\,
            I => dds_state_1
        );

    \I__11422\ : Odrv4
    port map (
            O => \N__50276\,
            I => dds_state_1
        );

    \I__11421\ : IoInMux
    port map (
            O => \N__50263\,
            I => \N__50260\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__50260\,
            I => \N__50257\
        );

    \I__11419\ : IoSpan4Mux
    port map (
            O => \N__50257\,
            I => \N__50254\
        );

    \I__11418\ : Sp12to4
    port map (
            O => \N__50254\,
            I => \N__50251\
        );

    \I__11417\ : Span12Mux_s6_v
    port map (
            O => \N__50251\,
            I => \N__50248\
        );

    \I__11416\ : Odrv12
    port map (
            O => \N__50248\,
            I => \DDS_CS\
        );

    \I__11415\ : CEMux
    port map (
            O => \N__50245\,
            I => \N__50242\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__50242\,
            I => \N__50239\
        );

    \I__11413\ : Span4Mux_v
    port map (
            O => \N__50239\,
            I => \N__50236\
        );

    \I__11412\ : Odrv4
    port map (
            O => \N__50236\,
            I => \SIG_DDS.n9_adj_1490\
        );

    \I__11411\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50230\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__50230\,
            I => \N__50227\
        );

    \I__11409\ : Span4Mux_v
    port map (
            O => \N__50227\,
            I => \N__50224\
        );

    \I__11408\ : Odrv4
    port map (
            O => \N__50224\,
            I => buf_data_iac_23
        );

    \I__11407\ : CascadeMux
    port map (
            O => \N__50221\,
            I => \N__50218\
        );

    \I__11406\ : InMux
    port map (
            O => \N__50218\,
            I => \N__50215\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__50215\,
            I => \N__50212\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__50212\,
            I => \N__50209\
        );

    \I__11403\ : Sp12to4
    port map (
            O => \N__50209\,
            I => \N__50206\
        );

    \I__11402\ : Span12Mux_v
    port map (
            O => \N__50206\,
            I => \N__50203\
        );

    \I__11401\ : Odrv12
    port map (
            O => \N__50203\,
            I => n22595
        );

    \I__11400\ : InMux
    port map (
            O => \N__50200\,
            I => \N__50195\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50199\,
            I => \N__50192\
        );

    \I__11398\ : InMux
    port map (
            O => \N__50198\,
            I => \N__50189\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__50195\,
            I => \N__50185\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__50192\,
            I => \N__50180\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__50189\,
            I => \N__50180\
        );

    \I__11394\ : InMux
    port map (
            O => \N__50188\,
            I => \N__50177\
        );

    \I__11393\ : Span4Mux_v
    port map (
            O => \N__50185\,
            I => \N__50174\
        );

    \I__11392\ : Span4Mux_v
    port map (
            O => \N__50180\,
            I => \N__50169\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__50177\,
            I => \N__50169\
        );

    \I__11390\ : Span4Mux_h
    port map (
            O => \N__50174\,
            I => \N__50165\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__50169\,
            I => \N__50162\
        );

    \I__11388\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50159\
        );

    \I__11387\ : Span4Mux_v
    port map (
            O => \N__50165\,
            I => \N__50156\
        );

    \I__11386\ : Span4Mux_v
    port map (
            O => \N__50162\,
            I => \N__50153\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__50159\,
            I => \N__50150\
        );

    \I__11384\ : Sp12to4
    port map (
            O => \N__50156\,
            I => \N__50143\
        );

    \I__11383\ : Sp12to4
    port map (
            O => \N__50153\,
            I => \N__50143\
        );

    \I__11382\ : Span12Mux_v
    port map (
            O => \N__50150\,
            I => \N__50143\
        );

    \I__11381\ : Odrv12
    port map (
            O => \N__50143\,
            I => \ICE_SPI_MOSI\
        );

    \I__11380\ : SRMux
    port map (
            O => \N__50140\,
            I => \N__50137\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__50137\,
            I => \N__50134\
        );

    \I__11378\ : Odrv4
    port map (
            O => \N__50134\,
            I => \comm_spi.imosi_N_840\
        );

    \I__11377\ : InMux
    port map (
            O => \N__50131\,
            I => n20630
        );

    \I__11376\ : InMux
    port map (
            O => \N__50128\,
            I => \N__50124\
        );

    \I__11375\ : CascadeMux
    port map (
            O => \N__50127\,
            I => \N__50121\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__50124\,
            I => \N__50118\
        );

    \I__11373\ : InMux
    port map (
            O => \N__50121\,
            I => \N__50114\
        );

    \I__11372\ : Span4Mux_v
    port map (
            O => \N__50118\,
            I => \N__50111\
        );

    \I__11371\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50108\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__50114\,
            I => \N__50105\
        );

    \I__11369\ : Span4Mux_h
    port map (
            O => \N__50111\,
            I => \N__50102\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__50108\,
            I => \N__50097\
        );

    \I__11367\ : Span4Mux_h
    port map (
            O => \N__50105\,
            I => \N__50097\
        );

    \I__11366\ : Odrv4
    port map (
            O => \N__50102\,
            I => data_cntvec_10
        );

    \I__11365\ : Odrv4
    port map (
            O => \N__50097\,
            I => data_cntvec_10
        );

    \I__11364\ : InMux
    port map (
            O => \N__50092\,
            I => n20631
        );

    \I__11363\ : InMux
    port map (
            O => \N__50089\,
            I => n20632
        );

    \I__11362\ : InMux
    port map (
            O => \N__50086\,
            I => \N__50083\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__50083\,
            I => \N__50079\
        );

    \I__11360\ : InMux
    port map (
            O => \N__50082\,
            I => \N__50076\
        );

    \I__11359\ : Span4Mux_h
    port map (
            O => \N__50079\,
            I => \N__50073\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__50076\,
            I => data_cntvec_12
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__50073\,
            I => data_cntvec_12
        );

    \I__11356\ : InMux
    port map (
            O => \N__50068\,
            I => n20633
        );

    \I__11355\ : InMux
    port map (
            O => \N__50065\,
            I => \N__50062\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__50062\,
            I => \N__50059\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__50059\,
            I => \N__50055\
        );

    \I__11352\ : InMux
    port map (
            O => \N__50058\,
            I => \N__50052\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__50055\,
            I => \N__50049\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__50052\,
            I => data_cntvec_13
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__50049\,
            I => data_cntvec_13
        );

    \I__11348\ : InMux
    port map (
            O => \N__50044\,
            I => n20634
        );

    \I__11347\ : InMux
    port map (
            O => \N__50041\,
            I => n20635
        );

    \I__11346\ : InMux
    port map (
            O => \N__50038\,
            I => n20636
        );

    \I__11345\ : InMux
    port map (
            O => \N__50035\,
            I => \N__50031\
        );

    \I__11344\ : InMux
    port map (
            O => \N__50034\,
            I => \N__50028\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__50031\,
            I => \N__50025\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__50028\,
            I => data_cntvec_15
        );

    \I__11341\ : Odrv4
    port map (
            O => \N__50025\,
            I => data_cntvec_15
        );

    \I__11340\ : InMux
    port map (
            O => \N__50020\,
            I => \N__50014\
        );

    \I__11339\ : CEMux
    port map (
            O => \N__50019\,
            I => \N__50010\
        );

    \I__11338\ : CEMux
    port map (
            O => \N__50018\,
            I => \N__50007\
        );

    \I__11337\ : CEMux
    port map (
            O => \N__50017\,
            I => \N__50004\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__50014\,
            I => \N__50001\
        );

    \I__11335\ : CEMux
    port map (
            O => \N__50013\,
            I => \N__49998\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__50010\,
            I => \N__49995\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__50007\,
            I => \N__49992\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__50004\,
            I => \N__49989\
        );

    \I__11331\ : Span4Mux_v
    port map (
            O => \N__50001\,
            I => \N__49986\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__49998\,
            I => \N__49983\
        );

    \I__11329\ : Span4Mux_h
    port map (
            O => \N__49995\,
            I => \N__49978\
        );

    \I__11328\ : Span4Mux_h
    port map (
            O => \N__49992\,
            I => \N__49978\
        );

    \I__11327\ : Span4Mux_v
    port map (
            O => \N__49989\,
            I => \N__49973\
        );

    \I__11326\ : Span4Mux_v
    port map (
            O => \N__49986\,
            I => \N__49973\
        );

    \I__11325\ : Span4Mux_h
    port map (
            O => \N__49983\,
            I => \N__49970\
        );

    \I__11324\ : Sp12to4
    port map (
            O => \N__49978\,
            I => \N__49967\
        );

    \I__11323\ : Span4Mux_h
    port map (
            O => \N__49973\,
            I => \N__49964\
        );

    \I__11322\ : Odrv4
    port map (
            O => \N__49970\,
            I => n12394
        );

    \I__11321\ : Odrv12
    port map (
            O => \N__49967\,
            I => n12394
        );

    \I__11320\ : Odrv4
    port map (
            O => \N__49964\,
            I => n12394
        );

    \I__11319\ : SRMux
    port map (
            O => \N__49957\,
            I => \N__49953\
        );

    \I__11318\ : SRMux
    port map (
            O => \N__49956\,
            I => \N__49950\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__49953\,
            I => \N__49947\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__49950\,
            I => \N__49944\
        );

    \I__11315\ : Span4Mux_v
    port map (
            O => \N__49947\,
            I => \N__49939\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__49944\,
            I => \N__49936\
        );

    \I__11313\ : SRMux
    port map (
            O => \N__49943\,
            I => \N__49933\
        );

    \I__11312\ : SRMux
    port map (
            O => \N__49942\,
            I => \N__49930\
        );

    \I__11311\ : Span4Mux_h
    port map (
            O => \N__49939\,
            I => \N__49925\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__49936\,
            I => \N__49925\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__49933\,
            I => \N__49922\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__49930\,
            I => \N__49919\
        );

    \I__11307\ : Span4Mux_h
    port map (
            O => \N__49925\,
            I => \N__49912\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__49922\,
            I => \N__49912\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__49919\,
            I => \N__49912\
        );

    \I__11304\ : Odrv4
    port map (
            O => \N__49912\,
            I => n15431
        );

    \I__11303\ : InMux
    port map (
            O => \N__49909\,
            I => \N__49906\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__49906\,
            I => \N__49903\
        );

    \I__11301\ : Span4Mux_h
    port map (
            O => \N__49903\,
            I => \N__49900\
        );

    \I__11300\ : Odrv4
    port map (
            O => \N__49900\,
            I => n23480
        );

    \I__11299\ : IoInMux
    port map (
            O => \N__49897\,
            I => \N__49894\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__49894\,
            I => \N__49891\
        );

    \I__11297\ : IoSpan4Mux
    port map (
            O => \N__49891\,
            I => \N__49888\
        );

    \I__11296\ : IoSpan4Mux
    port map (
            O => \N__49888\,
            I => \N__49885\
        );

    \I__11295\ : Span4Mux_s1_v
    port map (
            O => \N__49885\,
            I => \N__49881\
        );

    \I__11294\ : CascadeMux
    port map (
            O => \N__49884\,
            I => \N__49878\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__49881\,
            I => \N__49875\
        );

    \I__11292\ : InMux
    port map (
            O => \N__49878\,
            I => \N__49872\
        );

    \I__11291\ : Span4Mux_v
    port map (
            O => \N__49875\,
            I => \N__49867\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__49872\,
            I => \N__49867\
        );

    \I__11289\ : Span4Mux_h
    port map (
            O => \N__49867\,
            I => \N__49863\
        );

    \I__11288\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49860\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__49863\,
            I => \N__49857\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__49860\,
            I => \DDS_RNG_0\
        );

    \I__11285\ : Odrv4
    port map (
            O => \N__49857\,
            I => \DDS_RNG_0\
        );

    \I__11284\ : InMux
    port map (
            O => \N__49852\,
            I => \N__49849\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__49849\,
            I => \N__49845\
        );

    \I__11282\ : InMux
    port map (
            O => \N__49848\,
            I => \N__49841\
        );

    \I__11281\ : Span12Mux_h
    port map (
            O => \N__49845\,
            I => \N__49838\
        );

    \I__11280\ : InMux
    port map (
            O => \N__49844\,
            I => \N__49835\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__49841\,
            I => \acadc_skipCount_9\
        );

    \I__11278\ : Odrv12
    port map (
            O => \N__49838\,
            I => \acadc_skipCount_9\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__49835\,
            I => \acadc_skipCount_9\
        );

    \I__11276\ : CascadeMux
    port map (
            O => \N__49828\,
            I => \n22183_cascade_\
        );

    \I__11275\ : InMux
    port map (
            O => \N__49825\,
            I => n20622
        );

    \I__11274\ : InMux
    port map (
            O => \N__49822\,
            I => n20623
        );

    \I__11273\ : InMux
    port map (
            O => \N__49819\,
            I => \N__49816\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__49816\,
            I => \N__49812\
        );

    \I__11271\ : InMux
    port map (
            O => \N__49815\,
            I => \N__49808\
        );

    \I__11270\ : Span4Mux_h
    port map (
            O => \N__49812\,
            I => \N__49805\
        );

    \I__11269\ : InMux
    port map (
            O => \N__49811\,
            I => \N__49802\
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__49808\,
            I => data_cntvec_3
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__49805\,
            I => data_cntvec_3
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__49802\,
            I => data_cntvec_3
        );

    \I__11265\ : InMux
    port map (
            O => \N__49795\,
            I => n20624
        );

    \I__11264\ : InMux
    port map (
            O => \N__49792\,
            I => n20625
        );

    \I__11263\ : InMux
    port map (
            O => \N__49789\,
            I => n20626
        );

    \I__11262\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49783\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__49783\,
            I => \N__49779\
        );

    \I__11260\ : InMux
    port map (
            O => \N__49782\,
            I => \N__49775\
        );

    \I__11259\ : Span4Mux_h
    port map (
            O => \N__49779\,
            I => \N__49772\
        );

    \I__11258\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49769\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__49775\,
            I => data_cntvec_6
        );

    \I__11256\ : Odrv4
    port map (
            O => \N__49772\,
            I => data_cntvec_6
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__49769\,
            I => data_cntvec_6
        );

    \I__11254\ : InMux
    port map (
            O => \N__49762\,
            I => n20627
        );

    \I__11253\ : InMux
    port map (
            O => \N__49759\,
            I => n20628
        );

    \I__11252\ : InMux
    port map (
            O => \N__49756\,
            I => \N__49753\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__49753\,
            I => \N__49750\
        );

    \I__11250\ : Span4Mux_h
    port map (
            O => \N__49750\,
            I => \N__49747\
        );

    \I__11249\ : Span4Mux_h
    port map (
            O => \N__49747\,
            I => \N__49743\
        );

    \I__11248\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49739\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__49743\,
            I => \N__49736\
        );

    \I__11246\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49733\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__49739\,
            I => data_cntvec_8
        );

    \I__11244\ : Odrv4
    port map (
            O => \N__49736\,
            I => data_cntvec_8
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__49733\,
            I => data_cntvec_8
        );

    \I__11242\ : InMux
    port map (
            O => \N__49726\,
            I => \bfn_17_16_0_\
        );

    \I__11241\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49720\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49716\
        );

    \I__11239\ : InMux
    port map (
            O => \N__49719\,
            I => \N__49713\
        );

    \I__11238\ : Span4Mux_h
    port map (
            O => \N__49716\,
            I => \N__49710\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__49713\,
            I => data_idxvec_12
        );

    \I__11236\ : Odrv4
    port map (
            O => \N__49710\,
            I => data_idxvec_12
        );

    \I__11235\ : InMux
    port map (
            O => \N__49705\,
            I => \N__49702\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__49702\,
            I => \N__49699\
        );

    \I__11233\ : Span4Mux_v
    port map (
            O => \N__49699\,
            I => \N__49696\
        );

    \I__11232\ : Sp12to4
    port map (
            O => \N__49696\,
            I => \N__49693\
        );

    \I__11231\ : Odrv12
    port map (
            O => \N__49693\,
            I => n22499
        );

    \I__11230\ : InMux
    port map (
            O => \N__49690\,
            I => \N__49687\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__49687\,
            I => \N__49684\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__49684\,
            I => \N__49679\
        );

    \I__11227\ : InMux
    port map (
            O => \N__49683\,
            I => \N__49674\
        );

    \I__11226\ : InMux
    port map (
            O => \N__49682\,
            I => \N__49674\
        );

    \I__11225\ : Odrv4
    port map (
            O => \N__49679\,
            I => \acadc_skipCount_6\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__49674\,
            I => \acadc_skipCount_6\
        );

    \I__11223\ : CascadeMux
    port map (
            O => \N__49669\,
            I => \N__49666\
        );

    \I__11222\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49663\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__49663\,
            I => \N__49660\
        );

    \I__11220\ : Span4Mux_h
    port map (
            O => \N__49660\,
            I => \N__49657\
        );

    \I__11219\ : Sp12to4
    port map (
            O => \N__49657\,
            I => \N__49652\
        );

    \I__11218\ : InMux
    port map (
            O => \N__49656\,
            I => \N__49647\
        );

    \I__11217\ : InMux
    port map (
            O => \N__49655\,
            I => \N__49647\
        );

    \I__11216\ : Odrv12
    port map (
            O => \N__49652\,
            I => req_data_cnt_6
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__49647\,
            I => req_data_cnt_6
        );

    \I__11214\ : CascadeMux
    port map (
            O => \N__49642\,
            I => \n23519_cascade_\
        );

    \I__11213\ : InMux
    port map (
            O => \N__49639\,
            I => \N__49636\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__49636\,
            I => \N__49633\
        );

    \I__11211\ : Span4Mux_h
    port map (
            O => \N__49633\,
            I => \N__49630\
        );

    \I__11210\ : Odrv4
    port map (
            O => \N__49630\,
            I => n23291
        );

    \I__11209\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49624\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__49624\,
            I => \N__49621\
        );

    \I__11207\ : Odrv12
    port map (
            O => \N__49621\,
            I => n111_adj_1726
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__49618\,
            I => \n30_adj_1724_cascade_\
        );

    \I__11205\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49612\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__49612\,
            I => \comm_buf_1_7_N_559_6\
        );

    \I__11203\ : InMux
    port map (
            O => \N__49609\,
            I => \N__49606\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__49606\,
            I => \N__49602\
        );

    \I__11201\ : InMux
    port map (
            O => \N__49605\,
            I => \N__49599\
        );

    \I__11200\ : Span4Mux_v
    port map (
            O => \N__49602\,
            I => \N__49596\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__49599\,
            I => data_idxvec_6
        );

    \I__11198\ : Odrv4
    port map (
            O => \N__49596\,
            I => data_idxvec_6
        );

    \I__11197\ : CascadeMux
    port map (
            O => \N__49591\,
            I => \n26_adj_1723_cascade_\
        );

    \I__11196\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49585\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__49585\,
            I => n23516
        );

    \I__11194\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49579\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__49579\,
            I => n23303
        );

    \I__11192\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49573\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__49573\,
            I => n23555
        );

    \I__11190\ : InMux
    port map (
            O => \N__49570\,
            I => \N__49564\
        );

    \I__11189\ : InMux
    port map (
            O => \N__49569\,
            I => \N__49552\
        );

    \I__11188\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49552\
        );

    \I__11187\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49552\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__49564\,
            I => \N__49549\
        );

    \I__11185\ : InMux
    port map (
            O => \N__49563\,
            I => \N__49546\
        );

    \I__11184\ : InMux
    port map (
            O => \N__49562\,
            I => \N__49543\
        );

    \I__11183\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49538\
        );

    \I__11182\ : InMux
    port map (
            O => \N__49560\,
            I => \N__49538\
        );

    \I__11181\ : InMux
    port map (
            O => \N__49559\,
            I => \N__49534\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__49552\,
            I => \N__49531\
        );

    \I__11179\ : Span4Mux_v
    port map (
            O => \N__49549\,
            I => \N__49522\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49522\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__49543\,
            I => \N__49522\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49522\
        );

    \I__11175\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49519\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__49534\,
            I => \N__49515\
        );

    \I__11173\ : Span4Mux_v
    port map (
            O => \N__49531\,
            I => \N__49510\
        );

    \I__11172\ : Span4Mux_v
    port map (
            O => \N__49522\,
            I => \N__49510\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__49519\,
            I => \N__49507\
        );

    \I__11170\ : InMux
    port map (
            O => \N__49518\,
            I => \N__49504\
        );

    \I__11169\ : Span4Mux_h
    port map (
            O => \N__49515\,
            I => \N__49499\
        );

    \I__11168\ : Span4Mux_h
    port map (
            O => \N__49510\,
            I => \N__49494\
        );

    \I__11167\ : Span4Mux_v
    port map (
            O => \N__49507\,
            I => \N__49494\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__49504\,
            I => \N__49491\
        );

    \I__11165\ : InMux
    port map (
            O => \N__49503\,
            I => \N__49488\
        );

    \I__11164\ : InMux
    port map (
            O => \N__49502\,
            I => \N__49485\
        );

    \I__11163\ : Span4Mux_h
    port map (
            O => \N__49499\,
            I => \N__49482\
        );

    \I__11162\ : Span4Mux_h
    port map (
            O => \N__49494\,
            I => \N__49479\
        );

    \I__11161\ : Span12Mux_v
    port map (
            O => \N__49491\,
            I => \N__49474\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__49488\,
            I => \N__49474\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__49485\,
            I => \N__49471\
        );

    \I__11158\ : Odrv4
    port map (
            O => \N__49482\,
            I => n18363
        );

    \I__11157\ : Odrv4
    port map (
            O => \N__49479\,
            I => n18363
        );

    \I__11156\ : Odrv12
    port map (
            O => \N__49474\,
            I => n18363
        );

    \I__11155\ : Odrv12
    port map (
            O => \N__49471\,
            I => n18363
        );

    \I__11154\ : InMux
    port map (
            O => \N__49462\,
            I => \N__49459\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__49459\,
            I => \N__49454\
        );

    \I__11152\ : InMux
    port map (
            O => \N__49458\,
            I => \N__49451\
        );

    \I__11151\ : InMux
    port map (
            O => \N__49457\,
            I => \N__49448\
        );

    \I__11150\ : Span12Mux_s10_h
    port map (
            O => \N__49454\,
            I => \N__49443\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__49451\,
            I => \N__49443\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__49448\,
            I => buf_dds1_4
        );

    \I__11147\ : Odrv12
    port map (
            O => \N__49443\,
            I => buf_dds1_4
        );

    \I__11146\ : CascadeMux
    port map (
            O => \N__49438\,
            I => \N__49432\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__49437\,
            I => \N__49429\
        );

    \I__11144\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49424\
        );

    \I__11143\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49424\
        );

    \I__11142\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49421\
        );

    \I__11141\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49418\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__49424\,
            I => \N__49413\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__49421\,
            I => \N__49413\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__49418\,
            I => \N__49409\
        );

    \I__11137\ : Span12Mux_h
    port map (
            O => \N__49413\,
            I => \N__49406\
        );

    \I__11136\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49403\
        );

    \I__11135\ : Odrv4
    port map (
            O => \N__49409\,
            I => \iac_raw_buf_N_823\
        );

    \I__11134\ : Odrv12
    port map (
            O => \N__49406\,
            I => \iac_raw_buf_N_823\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49403\,
            I => \iac_raw_buf_N_823\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49396\,
            I => \N__49393\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__49393\,
            I => \N__49389\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49392\,
            I => \N__49385\
        );

    \I__11129\ : Span4Mux_h
    port map (
            O => \N__49389\,
            I => \N__49382\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49388\,
            I => \N__49379\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__49385\,
            I => data_cntvec_0
        );

    \I__11126\ : Odrv4
    port map (
            O => \N__49382\,
            I => data_cntvec_0
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__49379\,
            I => data_cntvec_0
        );

    \I__11124\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49369\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__49369\,
            I => n22351
        );

    \I__11122\ : CascadeMux
    port map (
            O => \N__49366\,
            I => \n4_adj_1709_cascade_\
        );

    \I__11121\ : CascadeMux
    port map (
            O => \N__49363\,
            I => \N__49359\
        );

    \I__11120\ : CascadeMux
    port map (
            O => \N__49362\,
            I => \N__49356\
        );

    \I__11119\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49351\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49351\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__49351\,
            I => n35
        );

    \I__11116\ : InMux
    port map (
            O => \N__49348\,
            I => \N__49345\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__49345\,
            I => n12_adj_1802
        );

    \I__11114\ : InMux
    port map (
            O => \N__49342\,
            I => \N__49339\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__49339\,
            I => \N__49336\
        );

    \I__11112\ : Span4Mux_h
    port map (
            O => \N__49336\,
            I => \N__49333\
        );

    \I__11111\ : Odrv4
    port map (
            O => \N__49333\,
            I => \comm_buf_1_7_N_559_3\
        );

    \I__11110\ : InMux
    port map (
            O => \N__49330\,
            I => \N__49327\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__49327\,
            I => \N__49323\
        );

    \I__11108\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49319\
        );

    \I__11107\ : Span4Mux_h
    port map (
            O => \N__49323\,
            I => \N__49315\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49312\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__49319\,
            I => \N__49308\
        );

    \I__11104\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49305\
        );

    \I__11103\ : Span4Mux_h
    port map (
            O => \N__49315\,
            I => \N__49300\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__49312\,
            I => \N__49300\
        );

    \I__11101\ : CascadeMux
    port map (
            O => \N__49311\,
            I => \N__49297\
        );

    \I__11100\ : Span4Mux_h
    port map (
            O => \N__49308\,
            I => \N__49294\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__49305\,
            I => \N__49289\
        );

    \I__11098\ : Span4Mux_v
    port map (
            O => \N__49300\,
            I => \N__49286\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49297\,
            I => \N__49283\
        );

    \I__11096\ : Span4Mux_v
    port map (
            O => \N__49294\,
            I => \N__49280\
        );

    \I__11095\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49277\
        );

    \I__11094\ : CascadeMux
    port map (
            O => \N__49292\,
            I => \N__49274\
        );

    \I__11093\ : Span4Mux_h
    port map (
            O => \N__49289\,
            I => \N__49268\
        );

    \I__11092\ : Span4Mux_h
    port map (
            O => \N__49286\,
            I => \N__49268\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__49283\,
            I => \N__49261\
        );

    \I__11090\ : Sp12to4
    port map (
            O => \N__49280\,
            I => \N__49261\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__49277\,
            I => \N__49261\
        );

    \I__11088\ : InMux
    port map (
            O => \N__49274\,
            I => \N__49258\
        );

    \I__11087\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49255\
        );

    \I__11086\ : Sp12to4
    port map (
            O => \N__49268\,
            I => \N__49250\
        );

    \I__11085\ : Span12Mux_v
    port map (
            O => \N__49261\,
            I => \N__49250\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__49258\,
            I => comm_buf_1_3
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__49255\,
            I => comm_buf_1_3
        );

    \I__11082\ : Odrv12
    port map (
            O => \N__49250\,
            I => comm_buf_1_3
        );

    \I__11081\ : CascadeMux
    port map (
            O => \N__49243\,
            I => \N__49240\
        );

    \I__11080\ : InMux
    port map (
            O => \N__49240\,
            I => \N__49236\
        );

    \I__11079\ : InMux
    port map (
            O => \N__49239\,
            I => \N__49233\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__49236\,
            I => \N__49225\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__49233\,
            I => \N__49225\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49232\,
            I => \N__49222\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49231\,
            I => \N__49218\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49230\,
            I => \N__49215\
        );

    \I__11073\ : Span4Mux_v
    port map (
            O => \N__49225\,
            I => \N__49211\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__49222\,
            I => \N__49208\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49221\,
            I => \N__49205\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__49218\,
            I => \N__49202\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__49215\,
            I => \N__49199\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49214\,
            I => \N__49196\
        );

    \I__11067\ : Span4Mux_v
    port map (
            O => \N__49211\,
            I => \N__49193\
        );

    \I__11066\ : Span4Mux_v
    port map (
            O => \N__49208\,
            I => \N__49188\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__49205\,
            I => \N__49188\
        );

    \I__11064\ : Span4Mux_h
    port map (
            O => \N__49202\,
            I => \N__49185\
        );

    \I__11063\ : Span4Mux_v
    port map (
            O => \N__49199\,
            I => \N__49182\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__49196\,
            I => \N__49179\
        );

    \I__11061\ : Sp12to4
    port map (
            O => \N__49193\,
            I => \N__49176\
        );

    \I__11060\ : Span4Mux_h
    port map (
            O => \N__49188\,
            I => \N__49173\
        );

    \I__11059\ : Span4Mux_h
    port map (
            O => \N__49185\,
            I => \N__49170\
        );

    \I__11058\ : Sp12to4
    port map (
            O => \N__49182\,
            I => \N__49165\
        );

    \I__11057\ : Span12Mux_h
    port map (
            O => \N__49179\,
            I => \N__49165\
        );

    \I__11056\ : Span12Mux_h
    port map (
            O => \N__49176\,
            I => \N__49162\
        );

    \I__11055\ : Span4Mux_v
    port map (
            O => \N__49173\,
            I => \N__49159\
        );

    \I__11054\ : Odrv4
    port map (
            O => \N__49170\,
            I => comm_buf_1_6
        );

    \I__11053\ : Odrv12
    port map (
            O => \N__49165\,
            I => comm_buf_1_6
        );

    \I__11052\ : Odrv12
    port map (
            O => \N__49162\,
            I => comm_buf_1_6
        );

    \I__11051\ : Odrv4
    port map (
            O => \N__49159\,
            I => comm_buf_1_6
        );

    \I__11050\ : CascadeMux
    port map (
            O => \N__49150\,
            I => \N__49147\
        );

    \I__11049\ : InMux
    port map (
            O => \N__49147\,
            I => \N__49143\
        );

    \I__11048\ : InMux
    port map (
            O => \N__49146\,
            I => \N__49137\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__49143\,
            I => \N__49134\
        );

    \I__11046\ : CascadeMux
    port map (
            O => \N__49142\,
            I => \N__49130\
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__49141\,
            I => \N__49126\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__49140\,
            I => \N__49123\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__49119\
        );

    \I__11042\ : Span4Mux_v
    port map (
            O => \N__49134\,
            I => \N__49116\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__49133\,
            I => \N__49113\
        );

    \I__11040\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49110\
        );

    \I__11039\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49107\
        );

    \I__11038\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49103\
        );

    \I__11037\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49100\
        );

    \I__11036\ : InMux
    port map (
            O => \N__49122\,
            I => \N__49097\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__49119\,
            I => \N__49094\
        );

    \I__11034\ : Span4Mux_v
    port map (
            O => \N__49116\,
            I => \N__49091\
        );

    \I__11033\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49088\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__49110\,
            I => \N__49082\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__49107\,
            I => \N__49082\
        );

    \I__11030\ : InMux
    port map (
            O => \N__49106\,
            I => \N__49079\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__49103\,
            I => \N__49076\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__49100\,
            I => \N__49073\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__49097\,
            I => \N__49066\
        );

    \I__11026\ : Span4Mux_v
    port map (
            O => \N__49094\,
            I => \N__49066\
        );

    \I__11025\ : Span4Mux_h
    port map (
            O => \N__49091\,
            I => \N__49066\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__49088\,
            I => \N__49063\
        );

    \I__11023\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49060\
        );

    \I__11022\ : Span4Mux_v
    port map (
            O => \N__49082\,
            I => \N__49057\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__49079\,
            I => \N__49052\
        );

    \I__11020\ : Span12Mux_v
    port map (
            O => \N__49076\,
            I => \N__49052\
        );

    \I__11019\ : Span4Mux_v
    port map (
            O => \N__49073\,
            I => \N__49047\
        );

    \I__11018\ : Span4Mux_h
    port map (
            O => \N__49066\,
            I => \N__49047\
        );

    \I__11017\ : Span12Mux_h
    port map (
            O => \N__49063\,
            I => \N__49042\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__49042\
        );

    \I__11015\ : Span4Mux_h
    port map (
            O => \N__49057\,
            I => \N__49039\
        );

    \I__11014\ : Odrv12
    port map (
            O => \N__49052\,
            I => comm_buf_1_0
        );

    \I__11013\ : Odrv4
    port map (
            O => \N__49047\,
            I => comm_buf_1_0
        );

    \I__11012\ : Odrv12
    port map (
            O => \N__49042\,
            I => comm_buf_1_0
        );

    \I__11011\ : Odrv4
    port map (
            O => \N__49039\,
            I => comm_buf_1_0
        );

    \I__11010\ : InMux
    port map (
            O => \N__49030\,
            I => \N__49027\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__49023\
        );

    \I__11008\ : InMux
    port map (
            O => \N__49026\,
            I => \N__49020\
        );

    \I__11007\ : Span4Mux_v
    port map (
            O => \N__49023\,
            I => \N__49017\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__49020\,
            I => data_idxvec_14
        );

    \I__11005\ : Odrv4
    port map (
            O => \N__49017\,
            I => data_idxvec_14
        );

    \I__11004\ : CascadeMux
    port map (
            O => \N__49012\,
            I => \N__49009\
        );

    \I__11003\ : InMux
    port map (
            O => \N__49009\,
            I => \N__49006\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__49006\,
            I => \N__49003\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__49003\,
            I => \N__49000\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__49000\,
            I => n22296
        );

    \I__10999\ : CascadeMux
    port map (
            O => \N__48997\,
            I => \n46_cascade_\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__48994\,
            I => \N__48990\
        );

    \I__10997\ : InMux
    port map (
            O => \N__48993\,
            I => \N__48987\
        );

    \I__10996\ : InMux
    port map (
            O => \N__48990\,
            I => \N__48983\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__48987\,
            I => \N__48980\
        );

    \I__10994\ : InMux
    port map (
            O => \N__48986\,
            I => \N__48977\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__48983\,
            I => \N__48974\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__48980\,
            I => \N__48971\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__48977\,
            I => comm_test_buf_24_0
        );

    \I__10990\ : Odrv12
    port map (
            O => \N__48974\,
            I => comm_test_buf_24_0
        );

    \I__10989\ : Odrv4
    port map (
            O => \N__48971\,
            I => comm_test_buf_24_0
        );

    \I__10988\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48961\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__48961\,
            I => \N__48958\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__48958\,
            I => \N__48954\
        );

    \I__10985\ : InMux
    port map (
            O => \N__48957\,
            I => \N__48951\
        );

    \I__10984\ : Span4Mux_h
    port map (
            O => \N__48954\,
            I => \N__48946\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__48951\,
            I => \N__48946\
        );

    \I__10982\ : Odrv4
    port map (
            O => \N__48946\,
            I => comm_test_buf_24_8
        );

    \I__10981\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48938\
        );

    \I__10980\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48935\
        );

    \I__10979\ : CascadeMux
    port map (
            O => \N__48941\,
            I => \N__48932\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__48938\,
            I => \N__48929\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__48935\,
            I => \N__48926\
        );

    \I__10976\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48923\
        );

    \I__10975\ : Span4Mux_v
    port map (
            O => \N__48929\,
            I => \N__48920\
        );

    \I__10974\ : Span4Mux_h
    port map (
            O => \N__48926\,
            I => \N__48917\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__48923\,
            I => \N__48912\
        );

    \I__10972\ : Span4Mux_h
    port map (
            O => \N__48920\,
            I => \N__48912\
        );

    \I__10971\ : Span4Mux_v
    port map (
            O => \N__48917\,
            I => \N__48909\
        );

    \I__10970\ : Span4Mux_h
    port map (
            O => \N__48912\,
            I => \N__48906\
        );

    \I__10969\ : Odrv4
    port map (
            O => \N__48909\,
            I => n14_adj_1662
        );

    \I__10968\ : Odrv4
    port map (
            O => \N__48906\,
            I => n14_adj_1662
        );

    \I__10967\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48897\
        );

    \I__10966\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48894\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__48897\,
            I => n4_adj_1749
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__48894\,
            I => n4_adj_1749
        );

    \I__10963\ : InMux
    port map (
            O => \N__48889\,
            I => \N__48886\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__48886\,
            I => \N__48883\
        );

    \I__10961\ : Odrv12
    port map (
            O => \N__48883\,
            I => n12_adj_1684
        );

    \I__10960\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48876\
        );

    \I__10959\ : InMux
    port map (
            O => \N__48879\,
            I => \N__48873\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__48876\,
            I => \N__48867\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__48873\,
            I => \N__48864\
        );

    \I__10956\ : InMux
    port map (
            O => \N__48872\,
            I => \N__48861\
        );

    \I__10955\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48858\
        );

    \I__10954\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48854\
        );

    \I__10953\ : Span4Mux_h
    port map (
            O => \N__48867\,
            I => \N__48849\
        );

    \I__10952\ : Span4Mux_v
    port map (
            O => \N__48864\,
            I => \N__48849\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__48861\,
            I => \N__48846\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__48858\,
            I => \N__48843\
        );

    \I__10949\ : InMux
    port map (
            O => \N__48857\,
            I => \N__48840\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__48854\,
            I => \N__48833\
        );

    \I__10947\ : Span4Mux_h
    port map (
            O => \N__48849\,
            I => \N__48833\
        );

    \I__10946\ : Span4Mux_h
    port map (
            O => \N__48846\,
            I => \N__48833\
        );

    \I__10945\ : Span4Mux_h
    port map (
            O => \N__48843\,
            I => \N__48830\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__48840\,
            I => \N__48827\
        );

    \I__10943\ : Span4Mux_v
    port map (
            O => \N__48833\,
            I => \N__48824\
        );

    \I__10942\ : Span4Mux_v
    port map (
            O => \N__48830\,
            I => \N__48821\
        );

    \I__10941\ : Odrv12
    port map (
            O => \N__48827\,
            I => n14_adj_1608
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__48824\,
            I => n14_adj_1608
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__48821\,
            I => n14_adj_1608
        );

    \I__10938\ : InMux
    port map (
            O => \N__48814\,
            I => \N__48811\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__48811\,
            I => \N__48804\
        );

    \I__10936\ : InMux
    port map (
            O => \N__48810\,
            I => \N__48801\
        );

    \I__10935\ : InMux
    port map (
            O => \N__48809\,
            I => \N__48791\
        );

    \I__10934\ : InMux
    port map (
            O => \N__48808\,
            I => \N__48791\
        );

    \I__10933\ : InMux
    port map (
            O => \N__48807\,
            I => \N__48791\
        );

    \I__10932\ : Span4Mux_v
    port map (
            O => \N__48804\,
            I => \N__48786\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__48801\,
            I => \N__48786\
        );

    \I__10930\ : InMux
    port map (
            O => \N__48800\,
            I => \N__48783\
        );

    \I__10929\ : InMux
    port map (
            O => \N__48799\,
            I => \N__48780\
        );

    \I__10928\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48777\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__48791\,
            I => \N__48774\
        );

    \I__10926\ : Span4Mux_v
    port map (
            O => \N__48786\,
            I => \N__48771\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__48783\,
            I => \N__48768\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__48780\,
            I => \N__48765\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__48777\,
            I => \N__48762\
        );

    \I__10922\ : Span4Mux_v
    port map (
            O => \N__48774\,
            I => \N__48759\
        );

    \I__10921\ : Span4Mux_v
    port map (
            O => \N__48771\,
            I => \N__48754\
        );

    \I__10920\ : Span4Mux_v
    port map (
            O => \N__48768\,
            I => \N__48754\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__48765\,
            I => \N__48751\
        );

    \I__10918\ : Span4Mux_v
    port map (
            O => \N__48762\,
            I => \N__48748\
        );

    \I__10917\ : Sp12to4
    port map (
            O => \N__48759\,
            I => \N__48745\
        );

    \I__10916\ : Sp12to4
    port map (
            O => \N__48754\,
            I => \N__48742\
        );

    \I__10915\ : Sp12to4
    port map (
            O => \N__48751\,
            I => \N__48739\
        );

    \I__10914\ : Sp12to4
    port map (
            O => \N__48748\,
            I => \N__48734\
        );

    \I__10913\ : Span12Mux_h
    port map (
            O => \N__48745\,
            I => \N__48734\
        );

    \I__10912\ : Span12Mux_h
    port map (
            O => \N__48742\,
            I => \N__48731\
        );

    \I__10911\ : Odrv12
    port map (
            O => \N__48739\,
            I => n13129
        );

    \I__10910\ : Odrv12
    port map (
            O => \N__48734\,
            I => n13129
        );

    \I__10909\ : Odrv12
    port map (
            O => \N__48731\,
            I => n13129
        );

    \I__10908\ : CascadeMux
    port map (
            O => \N__48724\,
            I => \N__48721\
        );

    \I__10907\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48716\
        );

    \I__10906\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48713\
        );

    \I__10905\ : InMux
    port map (
            O => \N__48719\,
            I => \N__48710\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__48716\,
            I => \N__48707\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__48713\,
            I => \N__48699\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__48710\,
            I => \N__48699\
        );

    \I__10901\ : Sp12to4
    port map (
            O => \N__48707\,
            I => \N__48699\
        );

    \I__10900\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48696\
        );

    \I__10899\ : Span12Mux_v
    port map (
            O => \N__48699\,
            I => \N__48693\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__48696\,
            I => \N__48689\
        );

    \I__10897\ : Span12Mux_h
    port map (
            O => \N__48693\,
            I => \N__48686\
        );

    \I__10896\ : InMux
    port map (
            O => \N__48692\,
            I => \N__48683\
        );

    \I__10895\ : Span4Mux_h
    port map (
            O => \N__48689\,
            I => \N__48680\
        );

    \I__10894\ : Odrv12
    port map (
            O => \N__48686\,
            I => \buf_cfgRTD_0\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__48683\,
            I => \buf_cfgRTD_0\
        );

    \I__10892\ : Odrv4
    port map (
            O => \N__48680\,
            I => \buf_cfgRTD_0\
        );

    \I__10891\ : CascadeMux
    port map (
            O => \N__48673\,
            I => \N__48670\
        );

    \I__10890\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48667\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__48667\,
            I => \N__48664\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__48664\,
            I => \N__48661\
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__48661\,
            I => n22238
        );

    \I__10886\ : CascadeMux
    port map (
            O => \N__48658\,
            I => \n22240_cascade_\
        );

    \I__10885\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48652\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__48652\,
            I => n23053
        );

    \I__10883\ : CascadeMux
    port map (
            O => \N__48649\,
            I => \n11280_cascade_\
        );

    \I__10882\ : CascadeMux
    port map (
            O => \N__48646\,
            I => \n12509_cascade_\
        );

    \I__10881\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48639\
        );

    \I__10880\ : InMux
    port map (
            O => \N__48642\,
            I => \N__48636\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__48639\,
            I => \N__48633\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__48636\,
            I => comm_length_2
        );

    \I__10877\ : Odrv4
    port map (
            O => \N__48633\,
            I => comm_length_2
        );

    \I__10876\ : CascadeMux
    port map (
            O => \N__48628\,
            I => \N__48625\
        );

    \I__10875\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48622\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__48622\,
            I => \N__48619\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__48619\,
            I => \N__48616\
        );

    \I__10872\ : Odrv4
    port map (
            O => \N__48616\,
            I => comm_length_0
        );

    \I__10871\ : InMux
    port map (
            O => \N__48613\,
            I => \N__48610\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__48610\,
            I => \N__48606\
        );

    \I__10869\ : InMux
    port map (
            O => \N__48609\,
            I => \N__48603\
        );

    \I__10868\ : Span4Mux_h
    port map (
            O => \N__48606\,
            I => \N__48597\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__48603\,
            I => \N__48597\
        );

    \I__10866\ : InMux
    port map (
            O => \N__48602\,
            I => \N__48594\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__48597\,
            I => \N__48591\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__48594\,
            I => buf_adcdata_vac_17
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__48591\,
            I => buf_adcdata_vac_17
        );

    \I__10862\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48583\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__48583\,
            I => \N__48580\
        );

    \I__10860\ : Span4Mux_h
    port map (
            O => \N__48580\,
            I => \N__48577\
        );

    \I__10859\ : Odrv4
    port map (
            O => \N__48577\,
            I => n23486
        );

    \I__10858\ : CascadeMux
    port map (
            O => \N__48574\,
            I => \N__48571\
        );

    \I__10857\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48568\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__48568\,
            I => \N__48565\
        );

    \I__10855\ : Span4Mux_v
    port map (
            O => \N__48565\,
            I => \N__48562\
        );

    \I__10854\ : Span4Mux_h
    port map (
            O => \N__48562\,
            I => \N__48558\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__48561\,
            I => \N__48555\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__48558\,
            I => \N__48552\
        );

    \I__10851\ : InMux
    port map (
            O => \N__48555\,
            I => \N__48549\
        );

    \I__10850\ : Odrv4
    port map (
            O => \N__48552\,
            I => buf_adcdata_vdc_17
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__48549\,
            I => buf_adcdata_vdc_17
        );

    \I__10848\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48523\
        );

    \I__10847\ : InMux
    port map (
            O => \N__48543\,
            I => \N__48523\
        );

    \I__10846\ : InMux
    port map (
            O => \N__48542\,
            I => \N__48523\
        );

    \I__10845\ : InMux
    port map (
            O => \N__48541\,
            I => \N__48523\
        );

    \I__10844\ : InMux
    port map (
            O => \N__48540\,
            I => \N__48514\
        );

    \I__10843\ : InMux
    port map (
            O => \N__48539\,
            I => \N__48514\
        );

    \I__10842\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48514\
        );

    \I__10841\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48514\
        );

    \I__10840\ : InMux
    port map (
            O => \N__48536\,
            I => \N__48493\
        );

    \I__10839\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48493\
        );

    \I__10838\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48493\
        );

    \I__10837\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48493\
        );

    \I__10836\ : InMux
    port map (
            O => \N__48532\,
            I => \N__48490\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__48523\,
            I => \N__48487\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__48514\,
            I => \N__48484\
        );

    \I__10833\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48475\
        );

    \I__10832\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48475\
        );

    \I__10831\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48475\
        );

    \I__10830\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48475\
        );

    \I__10829\ : InMux
    port map (
            O => \N__48509\,
            I => \N__48466\
        );

    \I__10828\ : InMux
    port map (
            O => \N__48508\,
            I => \N__48466\
        );

    \I__10827\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48466\
        );

    \I__10826\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48466\
        );

    \I__10825\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48457\
        );

    \I__10824\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48457\
        );

    \I__10823\ : InMux
    port map (
            O => \N__48503\,
            I => \N__48457\
        );

    \I__10822\ : InMux
    port map (
            O => \N__48502\,
            I => \N__48457\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__48493\,
            I => \N__48452\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__48490\,
            I => \N__48452\
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__48487\,
            I => n49
        );

    \I__10818\ : Odrv4
    port map (
            O => \N__48484\,
            I => n49
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__48475\,
            I => n49
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__48466\,
            I => n49
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__48457\,
            I => n49
        );

    \I__10814\ : Odrv4
    port map (
            O => \N__48452\,
            I => n49
        );

    \I__10813\ : InMux
    port map (
            O => \N__48439\,
            I => \bfn_17_8_0_\
        );

    \I__10812\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48432\
        );

    \I__10811\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48429\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__48432\,
            I => \N__48426\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__48429\,
            I => wdtick_cnt_24
        );

    \I__10808\ : Odrv4
    port map (
            O => \N__48426\,
            I => wdtick_cnt_24
        );

    \I__10807\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48418\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__48418\,
            I => \N__48397\
        );

    \I__10805\ : ClkMux
    port map (
            O => \N__48417\,
            I => \N__48352\
        );

    \I__10804\ : ClkMux
    port map (
            O => \N__48416\,
            I => \N__48352\
        );

    \I__10803\ : ClkMux
    port map (
            O => \N__48415\,
            I => \N__48352\
        );

    \I__10802\ : ClkMux
    port map (
            O => \N__48414\,
            I => \N__48352\
        );

    \I__10801\ : ClkMux
    port map (
            O => \N__48413\,
            I => \N__48352\
        );

    \I__10800\ : ClkMux
    port map (
            O => \N__48412\,
            I => \N__48352\
        );

    \I__10799\ : ClkMux
    port map (
            O => \N__48411\,
            I => \N__48352\
        );

    \I__10798\ : ClkMux
    port map (
            O => \N__48410\,
            I => \N__48352\
        );

    \I__10797\ : ClkMux
    port map (
            O => \N__48409\,
            I => \N__48352\
        );

    \I__10796\ : ClkMux
    port map (
            O => \N__48408\,
            I => \N__48352\
        );

    \I__10795\ : ClkMux
    port map (
            O => \N__48407\,
            I => \N__48352\
        );

    \I__10794\ : ClkMux
    port map (
            O => \N__48406\,
            I => \N__48352\
        );

    \I__10793\ : ClkMux
    port map (
            O => \N__48405\,
            I => \N__48352\
        );

    \I__10792\ : ClkMux
    port map (
            O => \N__48404\,
            I => \N__48352\
        );

    \I__10791\ : ClkMux
    port map (
            O => \N__48403\,
            I => \N__48352\
        );

    \I__10790\ : ClkMux
    port map (
            O => \N__48402\,
            I => \N__48352\
        );

    \I__10789\ : ClkMux
    port map (
            O => \N__48401\,
            I => \N__48352\
        );

    \I__10788\ : ClkMux
    port map (
            O => \N__48400\,
            I => \N__48352\
        );

    \I__10787\ : Glb2LocalMux
    port map (
            O => \N__48397\,
            I => \N__48352\
        );

    \I__10786\ : ClkMux
    port map (
            O => \N__48396\,
            I => \N__48352\
        );

    \I__10785\ : ClkMux
    port map (
            O => \N__48395\,
            I => \N__48352\
        );

    \I__10784\ : GlobalMux
    port map (
            O => \N__48352\,
            I => \DDS_MCLK1\
        );

    \I__10783\ : CEMux
    port map (
            O => \N__48349\,
            I => \N__48346\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__48346\,
            I => \N__48342\
        );

    \I__10781\ : CEMux
    port map (
            O => \N__48345\,
            I => \N__48339\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__48342\,
            I => \N__48332\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__48339\,
            I => \N__48332\
        );

    \I__10778\ : CEMux
    port map (
            O => \N__48338\,
            I => \N__48329\
        );

    \I__10777\ : CEMux
    port map (
            O => \N__48337\,
            I => \N__48326\
        );

    \I__10776\ : Span4Mux_v
    port map (
            O => \N__48332\,
            I => \N__48323\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__48329\,
            I => \N__48320\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__48326\,
            I => \N__48317\
        );

    \I__10773\ : Span4Mux_h
    port map (
            O => \N__48323\,
            I => \N__48314\
        );

    \I__10772\ : Span4Mux_h
    port map (
            O => \N__48320\,
            I => \N__48311\
        );

    \I__10771\ : Span4Mux_h
    port map (
            O => \N__48317\,
            I => \N__48308\
        );

    \I__10770\ : Odrv4
    port map (
            O => \N__48314\,
            I => n12366
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__48311\,
            I => n12366
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__48308\,
            I => n12366
        );

    \I__10767\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48298\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__48298\,
            I => n7_adj_1757
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__48295\,
            I => \n2562_cascade_\
        );

    \I__10764\ : SRMux
    port map (
            O => \N__48292\,
            I => \N__48288\
        );

    \I__10763\ : SRMux
    port map (
            O => \N__48291\,
            I => \N__48285\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__48288\,
            I => \N__48282\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__48285\,
            I => \N__48279\
        );

    \I__10760\ : Span4Mux_v
    port map (
            O => \N__48282\,
            I => \N__48276\
        );

    \I__10759\ : Odrv12
    port map (
            O => \N__48279\,
            I => n15378
        );

    \I__10758\ : Odrv4
    port map (
            O => \N__48276\,
            I => n15378
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__48271\,
            I => \N__48268\
        );

    \I__10756\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48265\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__48265\,
            I => n8_adj_1782
        );

    \I__10754\ : CEMux
    port map (
            O => \N__48262\,
            I => \N__48259\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48256\
        );

    \I__10752\ : Span4Mux_v
    port map (
            O => \N__48256\,
            I => \N__48253\
        );

    \I__10751\ : Odrv4
    port map (
            O => \N__48253\,
            I => n12540
        );

    \I__10750\ : InMux
    port map (
            O => \N__48250\,
            I => \N__48247\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48244\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__48244\,
            I => \N__48241\
        );

    \I__10747\ : Span4Mux_v
    port map (
            O => \N__48241\,
            I => \N__48238\
        );

    \I__10746\ : Odrv4
    port map (
            O => \N__48238\,
            I => n14_adj_1606
        );

    \I__10745\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48231\
        );

    \I__10744\ : InMux
    port map (
            O => \N__48234\,
            I => \N__48228\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__48231\,
            I => \N__48225\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__48228\,
            I => wdtick_cnt_16
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__48225\,
            I => wdtick_cnt_16
        );

    \I__10740\ : InMux
    port map (
            O => \N__48220\,
            I => \bfn_17_7_0_\
        );

    \I__10739\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48213\
        );

    \I__10738\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48210\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__48213\,
            I => wdtick_cnt_17
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48210\,
            I => wdtick_cnt_17
        );

    \I__10735\ : InMux
    port map (
            O => \N__48205\,
            I => n20782
        );

    \I__10734\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48198\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48195\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__48198\,
            I => \N__48192\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__48195\,
            I => wdtick_cnt_18
        );

    \I__10730\ : Odrv4
    port map (
            O => \N__48192\,
            I => wdtick_cnt_18
        );

    \I__10729\ : InMux
    port map (
            O => \N__48187\,
            I => n20783
        );

    \I__10728\ : CascadeMux
    port map (
            O => \N__48184\,
            I => \N__48180\
        );

    \I__10727\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48177\
        );

    \I__10726\ : InMux
    port map (
            O => \N__48180\,
            I => \N__48174\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__48177\,
            I => wdtick_cnt_19
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__48174\,
            I => wdtick_cnt_19
        );

    \I__10723\ : InMux
    port map (
            O => \N__48169\,
            I => n20784
        );

    \I__10722\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48162\
        );

    \I__10721\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48159\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__48162\,
            I => wdtick_cnt_20
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__48159\,
            I => wdtick_cnt_20
        );

    \I__10718\ : InMux
    port map (
            O => \N__48154\,
            I => n20785
        );

    \I__10717\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48147\
        );

    \I__10716\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48144\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__48147\,
            I => wdtick_cnt_21
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__48144\,
            I => wdtick_cnt_21
        );

    \I__10713\ : InMux
    port map (
            O => \N__48139\,
            I => n20786
        );

    \I__10712\ : InMux
    port map (
            O => \N__48136\,
            I => \N__48132\
        );

    \I__10711\ : InMux
    port map (
            O => \N__48135\,
            I => \N__48129\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__48132\,
            I => wdtick_cnt_22
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__48129\,
            I => wdtick_cnt_22
        );

    \I__10708\ : InMux
    port map (
            O => \N__48124\,
            I => n20787
        );

    \I__10707\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48117\
        );

    \I__10706\ : InMux
    port map (
            O => \N__48120\,
            I => \N__48114\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__48117\,
            I => wdtick_cnt_23
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__48114\,
            I => wdtick_cnt_23
        );

    \I__10703\ : InMux
    port map (
            O => \N__48109\,
            I => n20788
        );

    \I__10702\ : CascadeMux
    port map (
            O => \N__48106\,
            I => \N__48103\
        );

    \I__10701\ : InMux
    port map (
            O => \N__48103\,
            I => \N__48100\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__48100\,
            I => \N__48096\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48099\,
            I => \N__48093\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__48096\,
            I => wdtick_cnt_7
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__48093\,
            I => wdtick_cnt_7
        );

    \I__10696\ : InMux
    port map (
            O => \N__48088\,
            I => n20772
        );

    \I__10695\ : InMux
    port map (
            O => \N__48085\,
            I => \N__48081\
        );

    \I__10694\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48078\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48075\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__48078\,
            I => wdtick_cnt_8
        );

    \I__10691\ : Odrv4
    port map (
            O => \N__48075\,
            I => wdtick_cnt_8
        );

    \I__10690\ : InMux
    port map (
            O => \N__48070\,
            I => \bfn_17_6_0_\
        );

    \I__10689\ : InMux
    port map (
            O => \N__48067\,
            I => \N__48063\
        );

    \I__10688\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48060\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__48063\,
            I => wdtick_cnt_9
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__48060\,
            I => wdtick_cnt_9
        );

    \I__10685\ : InMux
    port map (
            O => \N__48055\,
            I => n20774
        );

    \I__10684\ : InMux
    port map (
            O => \N__48052\,
            I => \N__48048\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48051\,
            I => \N__48045\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__48048\,
            I => wdtick_cnt_10
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__48045\,
            I => wdtick_cnt_10
        );

    \I__10680\ : InMux
    port map (
            O => \N__48040\,
            I => n20775
        );

    \I__10679\ : InMux
    port map (
            O => \N__48037\,
            I => \N__48033\
        );

    \I__10678\ : InMux
    port map (
            O => \N__48036\,
            I => \N__48030\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__48033\,
            I => wdtick_cnt_11
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__48030\,
            I => wdtick_cnt_11
        );

    \I__10675\ : InMux
    port map (
            O => \N__48025\,
            I => n20776
        );

    \I__10674\ : InMux
    port map (
            O => \N__48022\,
            I => \N__48018\
        );

    \I__10673\ : InMux
    port map (
            O => \N__48021\,
            I => \N__48015\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__48018\,
            I => wdtick_cnt_12
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__48015\,
            I => wdtick_cnt_12
        );

    \I__10670\ : InMux
    port map (
            O => \N__48010\,
            I => n20777
        );

    \I__10669\ : InMux
    port map (
            O => \N__48007\,
            I => \N__48003\
        );

    \I__10668\ : InMux
    port map (
            O => \N__48006\,
            I => \N__48000\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__48003\,
            I => wdtick_cnt_13
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__48000\,
            I => wdtick_cnt_13
        );

    \I__10665\ : InMux
    port map (
            O => \N__47995\,
            I => n20778
        );

    \I__10664\ : InMux
    port map (
            O => \N__47992\,
            I => \N__47988\
        );

    \I__10663\ : InMux
    port map (
            O => \N__47991\,
            I => \N__47985\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__47988\,
            I => \N__47980\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__47985\,
            I => \N__47980\
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__47980\,
            I => wdtick_cnt_14
        );

    \I__10659\ : InMux
    port map (
            O => \N__47977\,
            I => n20779
        );

    \I__10658\ : InMux
    port map (
            O => \N__47974\,
            I => \N__47970\
        );

    \I__10657\ : InMux
    port map (
            O => \N__47973\,
            I => \N__47967\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__47970\,
            I => wdtick_cnt_15
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__47967\,
            I => wdtick_cnt_15
        );

    \I__10654\ : InMux
    port map (
            O => \N__47962\,
            I => n20780
        );

    \I__10653\ : InMux
    port map (
            O => \N__47959\,
            I => \N__47955\
        );

    \I__10652\ : InMux
    port map (
            O => \N__47958\,
            I => \N__47951\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__47955\,
            I => \N__47948\
        );

    \I__10650\ : InMux
    port map (
            O => \N__47954\,
            I => \N__47945\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__47951\,
            I => \comm_spi.n15330\
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__47948\,
            I => \comm_spi.n15330\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__47945\,
            I => \comm_spi.n15330\
        );

    \I__10646\ : InMux
    port map (
            O => \N__47938\,
            I => \N__47934\
        );

    \I__10645\ : InMux
    port map (
            O => \N__47937\,
            I => \N__47931\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__47934\,
            I => \N__47926\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__47931\,
            I => \N__47926\
        );

    \I__10642\ : Odrv4
    port map (
            O => \N__47926\,
            I => wdtick_cnt_0
        );

    \I__10641\ : InMux
    port map (
            O => \N__47923\,
            I => \bfn_17_5_0_\
        );

    \I__10640\ : InMux
    port map (
            O => \N__47920\,
            I => \N__47916\
        );

    \I__10639\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47913\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__47916\,
            I => wdtick_cnt_1
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__47913\,
            I => wdtick_cnt_1
        );

    \I__10636\ : InMux
    port map (
            O => \N__47908\,
            I => n20766
        );

    \I__10635\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47901\
        );

    \I__10634\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47898\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__47901\,
            I => wdtick_cnt_2
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__47898\,
            I => wdtick_cnt_2
        );

    \I__10631\ : InMux
    port map (
            O => \N__47893\,
            I => n20767
        );

    \I__10630\ : CascadeMux
    port map (
            O => \N__47890\,
            I => \N__47887\
        );

    \I__10629\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47884\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__47884\,
            I => \N__47880\
        );

    \I__10627\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47877\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__47880\,
            I => wdtick_cnt_3
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__47877\,
            I => wdtick_cnt_3
        );

    \I__10624\ : InMux
    port map (
            O => \N__47872\,
            I => n20768
        );

    \I__10623\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47865\
        );

    \I__10622\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47862\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__47865\,
            I => wdtick_cnt_4
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__47862\,
            I => wdtick_cnt_4
        );

    \I__10619\ : InMux
    port map (
            O => \N__47857\,
            I => n20769
        );

    \I__10618\ : CascadeMux
    port map (
            O => \N__47854\,
            I => \N__47851\
        );

    \I__10617\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47848\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__47848\,
            I => \N__47844\
        );

    \I__10615\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47841\
        );

    \I__10614\ : Odrv4
    port map (
            O => \N__47844\,
            I => wdtick_cnt_5
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__47841\,
            I => wdtick_cnt_5
        );

    \I__10612\ : InMux
    port map (
            O => \N__47836\,
            I => n20770
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__47833\,
            I => \N__47829\
        );

    \I__10610\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47826\
        );

    \I__10609\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47823\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__47826\,
            I => wdtick_cnt_6
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__47823\,
            I => wdtick_cnt_6
        );

    \I__10606\ : InMux
    port map (
            O => \N__47818\,
            I => n20771
        );

    \I__10605\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47810\
        );

    \I__10604\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47807\
        );

    \I__10603\ : InMux
    port map (
            O => \N__47813\,
            I => \N__47804\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__47810\,
            I => \N__47799\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__47807\,
            I => \N__47799\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__47804\,
            I => \N__47796\
        );

    \I__10599\ : Span4Mux_h
    port map (
            O => \N__47799\,
            I => \N__47793\
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__47796\,
            I => data_index_0
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__47793\,
            I => data_index_0
        );

    \I__10596\ : InMux
    port map (
            O => \N__47788\,
            I => \N__47785\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__47785\,
            I => \N__47780\
        );

    \I__10594\ : CascadeMux
    port map (
            O => \N__47784\,
            I => \N__47777\
        );

    \I__10593\ : CascadeMux
    port map (
            O => \N__47783\,
            I => \N__47766\
        );

    \I__10592\ : Span4Mux_v
    port map (
            O => \N__47780\,
            I => \N__47763\
        );

    \I__10591\ : InMux
    port map (
            O => \N__47777\,
            I => \N__47760\
        );

    \I__10590\ : CascadeMux
    port map (
            O => \N__47776\,
            I => \N__47757\
        );

    \I__10589\ : CascadeMux
    port map (
            O => \N__47775\,
            I => \N__47754\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__47774\,
            I => \N__47751\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__47773\,
            I => \N__47748\
        );

    \I__10586\ : CascadeMux
    port map (
            O => \N__47772\,
            I => \N__47745\
        );

    \I__10585\ : CascadeMux
    port map (
            O => \N__47771\,
            I => \N__47742\
        );

    \I__10584\ : CascadeMux
    port map (
            O => \N__47770\,
            I => \N__47739\
        );

    \I__10583\ : CascadeMux
    port map (
            O => \N__47769\,
            I => \N__47736\
        );

    \I__10582\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47733\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__47763\,
            I => \N__47728\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47728\
        );

    \I__10579\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47719\
        );

    \I__10578\ : InMux
    port map (
            O => \N__47754\,
            I => \N__47719\
        );

    \I__10577\ : InMux
    port map (
            O => \N__47751\,
            I => \N__47719\
        );

    \I__10576\ : InMux
    port map (
            O => \N__47748\,
            I => \N__47719\
        );

    \I__10575\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47710\
        );

    \I__10574\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47710\
        );

    \I__10573\ : InMux
    port map (
            O => \N__47739\,
            I => \N__47710\
        );

    \I__10572\ : InMux
    port map (
            O => \N__47736\,
            I => \N__47710\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__47733\,
            I => \N__47707\
        );

    \I__10570\ : Span4Mux_v
    port map (
            O => \N__47728\,
            I => \N__47704\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__47719\,
            I => \N__47699\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__47710\,
            I => \N__47699\
        );

    \I__10567\ : Odrv12
    port map (
            O => \N__47707\,
            I => n11254
        );

    \I__10566\ : Odrv4
    port map (
            O => \N__47704\,
            I => n11254
        );

    \I__10565\ : Odrv4
    port map (
            O => \N__47699\,
            I => n11254
        );

    \I__10564\ : CEMux
    port map (
            O => \N__47692\,
            I => \N__47688\
        );

    \I__10563\ : CEMux
    port map (
            O => \N__47691\,
            I => \N__47685\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__47688\,
            I => \N__47682\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__47685\,
            I => \N__47679\
        );

    \I__10560\ : Odrv12
    port map (
            O => \N__47682\,
            I => n13052
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__47679\,
            I => n13052
        );

    \I__10558\ : SRMux
    port map (
            O => \N__47674\,
            I => \N__47671\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__47671\,
            I => \N__47668\
        );

    \I__10556\ : Odrv4
    port map (
            O => \N__47668\,
            I => n15562
        );

    \I__10555\ : CascadeMux
    port map (
            O => \N__47665\,
            I => \n15562_cascade_\
        );

    \I__10554\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47656\
        );

    \I__10553\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47648\
        );

    \I__10552\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47648\
        );

    \I__10551\ : InMux
    port map (
            O => \N__47659\,
            I => \N__47648\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__47656\,
            I => \N__47645\
        );

    \I__10549\ : InMux
    port map (
            O => \N__47655\,
            I => \N__47642\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__47648\,
            I => \N__47637\
        );

    \I__10547\ : Span4Mux_h
    port map (
            O => \N__47645\,
            I => \N__47637\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__47642\,
            I => bit_cnt_0
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__47637\,
            I => bit_cnt_0
        );

    \I__10544\ : CEMux
    port map (
            O => \N__47632\,
            I => \N__47629\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__47629\,
            I => \N__47626\
        );

    \I__10542\ : Span4Mux_v
    port map (
            O => \N__47626\,
            I => \N__47622\
        );

    \I__10541\ : CEMux
    port map (
            O => \N__47625\,
            I => \N__47619\
        );

    \I__10540\ : Odrv4
    port map (
            O => \N__47622\,
            I => \SIG_DDS.n9\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__47619\,
            I => \SIG_DDS.n9\
        );

    \I__10538\ : IoInMux
    port map (
            O => \N__47614\,
            I => \N__47611\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__47611\,
            I => \N__47608\
        );

    \I__10536\ : Span4Mux_s2_v
    port map (
            O => \N__47608\,
            I => \N__47605\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__47605\,
            I => \N__47602\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__47602\,
            I => \N__47598\
        );

    \I__10533\ : CascadeMux
    port map (
            O => \N__47601\,
            I => \N__47595\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__47598\,
            I => \N__47592\
        );

    \I__10531\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47589\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__47592\,
            I => \DDS_SCK\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__47589\,
            I => \DDS_SCK\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__47584\,
            I => \N__47579\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__47583\,
            I => \N__47576\
        );

    \I__10526\ : CascadeMux
    port map (
            O => \N__47582\,
            I => \N__47572\
        );

    \I__10525\ : InMux
    port map (
            O => \N__47579\,
            I => \N__47569\
        );

    \I__10524\ : InMux
    port map (
            O => \N__47576\,
            I => \N__47566\
        );

    \I__10523\ : InMux
    port map (
            O => \N__47575\,
            I => \N__47563\
        );

    \I__10522\ : InMux
    port map (
            O => \N__47572\,
            I => \N__47560\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__47569\,
            I => \N__47555\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__47566\,
            I => \N__47555\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__47563\,
            I => \N__47550\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__47560\,
            I => \N__47550\
        );

    \I__10517\ : Span12Mux_h
    port map (
            O => \N__47555\,
            I => \N__47547\
        );

    \I__10516\ : Odrv12
    port map (
            O => \N__47550\,
            I => trig_dds0
        );

    \I__10515\ : Odrv12
    port map (
            O => \N__47547\,
            I => trig_dds0
        );

    \I__10514\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47538\
        );

    \I__10513\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47535\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__47538\,
            I => \comm_spi.imosi\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__47535\,
            I => \comm_spi.imosi\
        );

    \I__10510\ : SRMux
    port map (
            O => \N__47530\,
            I => \N__47527\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__47527\,
            I => \N__47524\
        );

    \I__10508\ : Odrv4
    port map (
            O => \N__47524\,
            I => \comm_spi.DOUT_7__N_834\
        );

    \I__10507\ : InMux
    port map (
            O => \N__47521\,
            I => \N__47518\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__47518\,
            I => \N__47512\
        );

    \I__10505\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47509\
        );

    \I__10504\ : InMux
    port map (
            O => \N__47516\,
            I => \N__47506\
        );

    \I__10503\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47503\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__47512\,
            I => \N__47498\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__47509\,
            I => \N__47498\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__47506\,
            I => \N__47495\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__47503\,
            I => \N__47492\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__47498\,
            I => \N__47489\
        );

    \I__10497\ : Span4Mux_h
    port map (
            O => \N__47495\,
            I => \N__47486\
        );

    \I__10496\ : Odrv12
    port map (
            O => \N__47492\,
            I => n14_adj_1609
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__47489\,
            I => n14_adj_1609
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__47486\,
            I => n14_adj_1609
        );

    \I__10493\ : InMux
    port map (
            O => \N__47479\,
            I => n20667
        );

    \I__10492\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47472\
        );

    \I__10491\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47469\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__47472\,
            I => \N__47466\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__47469\,
            I => data_idxvec_8
        );

    \I__10488\ : Odrv4
    port map (
            O => \N__47466\,
            I => data_idxvec_8
        );

    \I__10487\ : InMux
    port map (
            O => \N__47461\,
            I => \bfn_16_17_0_\
        );

    \I__10486\ : InMux
    port map (
            O => \N__47458\,
            I => n20669
        );

    \I__10485\ : InMux
    port map (
            O => \N__47455\,
            I => \N__47446\
        );

    \I__10484\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47446\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__47453\,
            I => \N__47443\
        );

    \I__10482\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47440\
        );

    \I__10481\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47437\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__47446\,
            I => \N__47434\
        );

    \I__10479\ : InMux
    port map (
            O => \N__47443\,
            I => \N__47431\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__47440\,
            I => \N__47428\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__47437\,
            I => \N__47425\
        );

    \I__10476\ : Span4Mux_h
    port map (
            O => \N__47434\,
            I => \N__47419\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__47431\,
            I => \N__47419\
        );

    \I__10474\ : Span4Mux_v
    port map (
            O => \N__47428\,
            I => \N__47416\
        );

    \I__10473\ : Span4Mux_v
    port map (
            O => \N__47425\,
            I => \N__47413\
        );

    \I__10472\ : InMux
    port map (
            O => \N__47424\,
            I => \N__47410\
        );

    \I__10471\ : Span4Mux_v
    port map (
            O => \N__47419\,
            I => \N__47407\
        );

    \I__10470\ : Span4Mux_h
    port map (
            O => \N__47416\,
            I => \N__47402\
        );

    \I__10469\ : Span4Mux_v
    port map (
            O => \N__47413\,
            I => \N__47402\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__47410\,
            I => \N__47397\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__47407\,
            I => \N__47397\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__47402\,
            I => n14_adj_1655
        );

    \I__10465\ : Odrv4
    port map (
            O => \N__47397\,
            I => n14_adj_1655
        );

    \I__10464\ : InMux
    port map (
            O => \N__47392\,
            I => \N__47388\
        );

    \I__10463\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47385\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__47388\,
            I => data_idxvec_10
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__47385\,
            I => data_idxvec_10
        );

    \I__10460\ : InMux
    port map (
            O => \N__47380\,
            I => n20670
        );

    \I__10459\ : InMux
    port map (
            O => \N__47377\,
            I => n20671
        );

    \I__10458\ : InMux
    port map (
            O => \N__47374\,
            I => \N__47368\
        );

    \I__10457\ : InMux
    port map (
            O => \N__47373\,
            I => \N__47368\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47364\
        );

    \I__10455\ : InMux
    port map (
            O => \N__47367\,
            I => \N__47360\
        );

    \I__10454\ : Span4Mux_v
    port map (
            O => \N__47364\,
            I => \N__47357\
        );

    \I__10453\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47353\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__47360\,
            I => \N__47349\
        );

    \I__10451\ : Span4Mux_v
    port map (
            O => \N__47357\,
            I => \N__47346\
        );

    \I__10450\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47343\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__47353\,
            I => \N__47340\
        );

    \I__10448\ : InMux
    port map (
            O => \N__47352\,
            I => \N__47337\
        );

    \I__10447\ : Span4Mux_h
    port map (
            O => \N__47349\,
            I => \N__47334\
        );

    \I__10446\ : Sp12to4
    port map (
            O => \N__47346\,
            I => \N__47329\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__47343\,
            I => \N__47329\
        );

    \I__10444\ : Span4Mux_h
    port map (
            O => \N__47340\,
            I => \N__47324\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__47337\,
            I => \N__47324\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__47334\,
            I => n14_adj_1653
        );

    \I__10441\ : Odrv12
    port map (
            O => \N__47329\,
            I => n14_adj_1653
        );

    \I__10440\ : Odrv4
    port map (
            O => \N__47324\,
            I => n14_adj_1653
        );

    \I__10439\ : InMux
    port map (
            O => \N__47317\,
            I => n20672
        );

    \I__10438\ : InMux
    port map (
            O => \N__47314\,
            I => n20673
        );

    \I__10437\ : InMux
    port map (
            O => \N__47311\,
            I => n20674
        );

    \I__10436\ : InMux
    port map (
            O => \N__47308\,
            I => \N__47305\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__47305\,
            I => \N__47302\
        );

    \I__10434\ : Span4Mux_v
    port map (
            O => \N__47302\,
            I => \N__47299\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__47299\,
            I => n14_adj_1607
        );

    \I__10432\ : InMux
    port map (
            O => \N__47296\,
            I => n20675
        );

    \I__10431\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47290\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__47290\,
            I => \N__47286\
        );

    \I__10429\ : CascadeMux
    port map (
            O => \N__47289\,
            I => \N__47283\
        );

    \I__10428\ : Span4Mux_h
    port map (
            O => \N__47286\,
            I => \N__47280\
        );

    \I__10427\ : InMux
    port map (
            O => \N__47283\,
            I => \N__47277\
        );

    \I__10426\ : Span4Mux_h
    port map (
            O => \N__47280\,
            I => \N__47274\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__47277\,
            I => data_idxvec_15
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__47274\,
            I => data_idxvec_15
        );

    \I__10423\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47264\
        );

    \I__10422\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47261\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__47267\,
            I => \N__47258\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__47261\,
            I => \N__47252\
        );

    \I__10418\ : InMux
    port map (
            O => \N__47258\,
            I => \N__47249\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__47255\,
            I => \N__47246\
        );

    \I__10416\ : Span4Mux_h
    port map (
            O => \N__47252\,
            I => \N__47243\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__47249\,
            I => \N__47236\
        );

    \I__10414\ : Span4Mux_h
    port map (
            O => \N__47246\,
            I => \N__47236\
        );

    \I__10413\ : Span4Mux_h
    port map (
            O => \N__47243\,
            I => \N__47236\
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__47236\,
            I => buf_dds0_4
        );

    \I__10411\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47229\
        );

    \I__10410\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47226\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47223\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__47226\,
            I => \N__47220\
        );

    \I__10407\ : Span4Mux_v
    port map (
            O => \N__47223\,
            I => \N__47214\
        );

    \I__10406\ : Span4Mux_h
    port map (
            O => \N__47220\,
            I => \N__47214\
        );

    \I__10405\ : InMux
    port map (
            O => \N__47219\,
            I => \N__47211\
        );

    \I__10404\ : Span4Mux_h
    port map (
            O => \N__47214\,
            I => \N__47208\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__47211\,
            I => buf_dds0_0
        );

    \I__10402\ : Odrv4
    port map (
            O => \N__47208\,
            I => buf_dds0_0
        );

    \I__10401\ : InMux
    port map (
            O => \N__47203\,
            I => \N__47199\
        );

    \I__10400\ : InMux
    port map (
            O => \N__47202\,
            I => \N__47196\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__47199\,
            I => \N__47193\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__47196\,
            I => data_idxvec_0
        );

    \I__10397\ : Odrv4
    port map (
            O => \N__47193\,
            I => data_idxvec_0
        );

    \I__10396\ : InMux
    port map (
            O => \N__47188\,
            I => \bfn_16_16_0_\
        );

    \I__10395\ : InMux
    port map (
            O => \N__47185\,
            I => \N__47182\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__47182\,
            I => \N__47179\
        );

    \I__10393\ : Span4Mux_v
    port map (
            O => \N__47179\,
            I => \N__47176\
        );

    \I__10392\ : Span4Mux_v
    port map (
            O => \N__47176\,
            I => \N__47172\
        );

    \I__10391\ : InMux
    port map (
            O => \N__47175\,
            I => \N__47169\
        );

    \I__10390\ : Sp12to4
    port map (
            O => \N__47172\,
            I => \N__47164\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__47169\,
            I => \N__47164\
        );

    \I__10388\ : Odrv12
    port map (
            O => \N__47164\,
            I => n14_adj_1613
        );

    \I__10387\ : InMux
    port map (
            O => \N__47161\,
            I => n20661
        );

    \I__10386\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47155\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__47155\,
            I => \N__47151\
        );

    \I__10384\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47148\
        );

    \I__10383\ : Span4Mux_v
    port map (
            O => \N__47151\,
            I => \N__47145\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__47148\,
            I => n14_adj_1612
        );

    \I__10381\ : Odrv4
    port map (
            O => \N__47145\,
            I => n14_adj_1612
        );

    \I__10380\ : InMux
    port map (
            O => \N__47140\,
            I => n20662
        );

    \I__10379\ : CascadeMux
    port map (
            O => \N__47137\,
            I => \N__47134\
        );

    \I__10378\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47130\
        );

    \I__10377\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47127\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__47130\,
            I => \N__47124\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__47127\,
            I => data_idxvec_3
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__47124\,
            I => data_idxvec_3
        );

    \I__10373\ : InMux
    port map (
            O => \N__47119\,
            I => n20663
        );

    \I__10372\ : InMux
    port map (
            O => \N__47116\,
            I => n20664
        );

    \I__10371\ : CascadeMux
    port map (
            O => \N__47113\,
            I => \N__47109\
        );

    \I__10370\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47106\
        );

    \I__10369\ : InMux
    port map (
            O => \N__47109\,
            I => \N__47103\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__47106\,
            I => \N__47100\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__47103\,
            I => \N__47094\
        );

    \I__10366\ : Span4Mux_h
    port map (
            O => \N__47100\,
            I => \N__47094\
        );

    \I__10365\ : InMux
    port map (
            O => \N__47099\,
            I => \N__47091\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__47094\,
            I => \N__47088\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__47091\,
            I => \N__47085\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__47088\,
            I => n14_adj_1661
        );

    \I__10361\ : Odrv12
    port map (
            O => \N__47085\,
            I => n14_adj_1661
        );

    \I__10360\ : InMux
    port map (
            O => \N__47080\,
            I => n20665
        );

    \I__10359\ : InMux
    port map (
            O => \N__47077\,
            I => \N__47073\
        );

    \I__10358\ : CascadeMux
    port map (
            O => \N__47076\,
            I => \N__47070\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__47073\,
            I => \N__47066\
        );

    \I__10356\ : InMux
    port map (
            O => \N__47070\,
            I => \N__47063\
        );

    \I__10355\ : InMux
    port map (
            O => \N__47069\,
            I => \N__47060\
        );

    \I__10354\ : Span4Mux_v
    port map (
            O => \N__47066\,
            I => \N__47057\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__47063\,
            I => \N__47052\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__47060\,
            I => \N__47052\
        );

    \I__10351\ : Span4Mux_h
    port map (
            O => \N__47057\,
            I => \N__47047\
        );

    \I__10350\ : Span4Mux_v
    port map (
            O => \N__47052\,
            I => \N__47047\
        );

    \I__10349\ : Odrv4
    port map (
            O => \N__47047\,
            I => n14_adj_1610
        );

    \I__10348\ : InMux
    port map (
            O => \N__47044\,
            I => n20666
        );

    \I__10347\ : CascadeMux
    port map (
            O => \N__47041\,
            I => \n26_adj_1580_cascade_\
        );

    \I__10346\ : InMux
    port map (
            O => \N__47038\,
            I => \N__47035\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__47035\,
            I => \N__47032\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__47032\,
            I => \N__47027\
        );

    \I__10343\ : InMux
    port map (
            O => \N__47031\,
            I => \N__47022\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47030\,
            I => \N__47022\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__47027\,
            I => \acadc_skipCount_0\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47022\,
            I => \acadc_skipCount_0\
        );

    \I__10339\ : CascadeMux
    port map (
            O => \N__47017\,
            I => \n23552_cascade_\
        );

    \I__10338\ : InMux
    port map (
            O => \N__47014\,
            I => \N__47010\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__47013\,
            I => \N__47006\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__47010\,
            I => \N__47003\
        );

    \I__10335\ : InMux
    port map (
            O => \N__47009\,
            I => \N__47000\
        );

    \I__10334\ : InMux
    port map (
            O => \N__47006\,
            I => \N__46997\
        );

    \I__10333\ : Odrv4
    port map (
            O => \N__47003\,
            I => req_data_cnt_0
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__47000\,
            I => req_data_cnt_0
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__46997\,
            I => req_data_cnt_0
        );

    \I__10330\ : InMux
    port map (
            O => \N__46990\,
            I => \N__46987\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__46987\,
            I => \N__46984\
        );

    \I__10328\ : Span4Mux_h
    port map (
            O => \N__46984\,
            I => \N__46981\
        );

    \I__10327\ : Span4Mux_h
    port map (
            O => \N__46981\,
            I => \N__46978\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__46978\,
            I => n16
        );

    \I__10325\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46972\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__46972\,
            I => \N__46969\
        );

    \I__10323\ : Span4Mux_v
    port map (
            O => \N__46969\,
            I => \N__46966\
        );

    \I__10322\ : Sp12to4
    port map (
            O => \N__46966\,
            I => \N__46963\
        );

    \I__10321\ : Odrv12
    port map (
            O => \N__46963\,
            I => n23300
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__46960\,
            I => \N__46957\
        );

    \I__10319\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46953\
        );

    \I__10318\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46950\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__46953\,
            I => \N__46947\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46943\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__46947\,
            I => \N__46940\
        );

    \I__10314\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46937\
        );

    \I__10313\ : Span12Mux_s9_v
    port map (
            O => \N__46943\,
            I => \N__46934\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__46940\,
            I => \N__46931\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__46937\,
            I => buf_adcdata_iac_8
        );

    \I__10310\ : Odrv12
    port map (
            O => \N__46934\,
            I => buf_adcdata_iac_8
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__46931\,
            I => buf_adcdata_iac_8
        );

    \I__10308\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46921\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__46921\,
            I => \N__46917\
        );

    \I__10306\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46914\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__46917\,
            I => \N__46911\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__46914\,
            I => \N__46907\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__46911\,
            I => \N__46904\
        );

    \I__10302\ : CascadeMux
    port map (
            O => \N__46910\,
            I => \N__46901\
        );

    \I__10301\ : Span4Mux_h
    port map (
            O => \N__46907\,
            I => \N__46898\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__46904\,
            I => \N__46895\
        );

    \I__10299\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46892\
        );

    \I__10298\ : Span4Mux_h
    port map (
            O => \N__46898\,
            I => \N__46889\
        );

    \I__10297\ : Span4Mux_h
    port map (
            O => \N__46895\,
            I => \N__46886\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__46892\,
            I => buf_adcdata_iac_15
        );

    \I__10295\ : Odrv4
    port map (
            O => \N__46889\,
            I => buf_adcdata_iac_15
        );

    \I__10294\ : Odrv4
    port map (
            O => \N__46886\,
            I => buf_adcdata_iac_15
        );

    \I__10293\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46876\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__46876\,
            I => \N__46873\
        );

    \I__10291\ : Span4Mux_h
    port map (
            O => \N__46873\,
            I => \N__46870\
        );

    \I__10290\ : Span4Mux_h
    port map (
            O => \N__46870\,
            I => \N__46867\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__46867\,
            I => n16_adj_1713
        );

    \I__10288\ : InMux
    port map (
            O => \N__46864\,
            I => \N__46861\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46858\
        );

    \I__10286\ : Span4Mux_v
    port map (
            O => \N__46858\,
            I => \N__46855\
        );

    \I__10285\ : Odrv4
    port map (
            O => \N__46855\,
            I => n22268
        );

    \I__10284\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46839\
        );

    \I__10283\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46836\
        );

    \I__10282\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46831\
        );

    \I__10281\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46831\
        );

    \I__10280\ : InMux
    port map (
            O => \N__46848\,
            I => \N__46826\
        );

    \I__10279\ : InMux
    port map (
            O => \N__46847\,
            I => \N__46826\
        );

    \I__10278\ : InMux
    port map (
            O => \N__46846\,
            I => \N__46821\
        );

    \I__10277\ : InMux
    port map (
            O => \N__46845\,
            I => \N__46821\
        );

    \I__10276\ : CascadeMux
    port map (
            O => \N__46844\,
            I => \N__46814\
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__46843\,
            I => \N__46811\
        );

    \I__10274\ : InMux
    port map (
            O => \N__46842\,
            I => \N__46807\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__46839\,
            I => \N__46804\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__46836\,
            I => \N__46799\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__46831\,
            I => \N__46799\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__46826\,
            I => \N__46794\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__46821\,
            I => \N__46794\
        );

    \I__10268\ : InMux
    port map (
            O => \N__46820\,
            I => \N__46791\
        );

    \I__10267\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46788\
        );

    \I__10266\ : InMux
    port map (
            O => \N__46818\,
            I => \N__46785\
        );

    \I__10265\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46782\
        );

    \I__10264\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46775\
        );

    \I__10263\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46775\
        );

    \I__10262\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46775\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__46807\,
            I => \N__46768\
        );

    \I__10260\ : Span4Mux_v
    port map (
            O => \N__46804\,
            I => \N__46768\
        );

    \I__10259\ : Span4Mux_v
    port map (
            O => \N__46799\,
            I => \N__46768\
        );

    \I__10258\ : Span4Mux_h
    port map (
            O => \N__46794\,
            I => \N__46765\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__46791\,
            I => n13141
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__46788\,
            I => n13141
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__46785\,
            I => n13141
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__46782\,
            I => n13141
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__46775\,
            I => n13141
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__46768\,
            I => n13141
        );

    \I__10251\ : Odrv4
    port map (
            O => \N__46765\,
            I => n13141
        );

    \I__10250\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46745\
        );

    \I__10249\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46742\
        );

    \I__10248\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46739\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__46745\,
            I => \N__46733\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46730\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__46739\,
            I => \N__46727\
        );

    \I__10244\ : InMux
    port map (
            O => \N__46738\,
            I => \N__46720\
        );

    \I__10243\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46720\
        );

    \I__10242\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46720\
        );

    \I__10241\ : Span4Mux_v
    port map (
            O => \N__46733\,
            I => \N__46717\
        );

    \I__10240\ : Span4Mux_v
    port map (
            O => \N__46730\,
            I => \N__46712\
        );

    \I__10239\ : Span4Mux_v
    port map (
            O => \N__46727\,
            I => \N__46712\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46709\
        );

    \I__10237\ : Span4Mux_v
    port map (
            O => \N__46717\,
            I => \N__46706\
        );

    \I__10236\ : Span4Mux_h
    port map (
            O => \N__46712\,
            I => \N__46701\
        );

    \I__10235\ : Span4Mux_v
    port map (
            O => \N__46709\,
            I => \N__46701\
        );

    \I__10234\ : Span4Mux_v
    port map (
            O => \N__46706\,
            I => \N__46698\
        );

    \I__10233\ : Sp12to4
    port map (
            O => \N__46701\,
            I => \N__46695\
        );

    \I__10232\ : Odrv4
    port map (
            O => \N__46698\,
            I => n12610
        );

    \I__10231\ : Odrv12
    port map (
            O => \N__46695\,
            I => n12610
        );

    \I__10230\ : CascadeMux
    port map (
            O => \N__46690\,
            I => \n12021_cascade_\
        );

    \I__10229\ : CEMux
    port map (
            O => \N__46687\,
            I => \N__46684\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__46684\,
            I => n12614
        );

    \I__10227\ : CascadeMux
    port map (
            O => \N__46681\,
            I => \n25_cascade_\
        );

    \I__10226\ : CEMux
    port map (
            O => \N__46678\,
            I => \N__46675\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46672\
        );

    \I__10224\ : Span4Mux_v
    port map (
            O => \N__46672\,
            I => \N__46669\
        );

    \I__10223\ : Sp12to4
    port map (
            O => \N__46669\,
            I => \N__46666\
        );

    \I__10222\ : Odrv12
    port map (
            O => \N__46666\,
            I => n12548
        );

    \I__10221\ : CascadeMux
    port map (
            O => \N__46663\,
            I => \N__46659\
        );

    \I__10220\ : CascadeMux
    port map (
            O => \N__46662\,
            I => \N__46655\
        );

    \I__10219\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46651\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__46658\,
            I => \N__46648\
        );

    \I__10217\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46643\
        );

    \I__10216\ : CascadeMux
    port map (
            O => \N__46654\,
            I => \N__46639\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__46651\,
            I => \N__46636\
        );

    \I__10214\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46633\
        );

    \I__10213\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46630\
        );

    \I__10212\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46626\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__46643\,
            I => \N__46623\
        );

    \I__10210\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46617\
        );

    \I__10209\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46614\
        );

    \I__10208\ : Span4Mux_v
    port map (
            O => \N__46636\,
            I => \N__46611\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__46633\,
            I => \N__46608\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__46630\,
            I => \N__46605\
        );

    \I__10205\ : CascadeMux
    port map (
            O => \N__46629\,
            I => \N__46602\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__46626\,
            I => \N__46599\
        );

    \I__10203\ : Span4Mux_v
    port map (
            O => \N__46623\,
            I => \N__46596\
        );

    \I__10202\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46593\
        );

    \I__10201\ : InMux
    port map (
            O => \N__46621\,
            I => \N__46588\
        );

    \I__10200\ : InMux
    port map (
            O => \N__46620\,
            I => \N__46588\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46585\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__46614\,
            I => \N__46582\
        );

    \I__10197\ : Span4Mux_h
    port map (
            O => \N__46611\,
            I => \N__46575\
        );

    \I__10196\ : Span4Mux_h
    port map (
            O => \N__46608\,
            I => \N__46575\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__46605\,
            I => \N__46575\
        );

    \I__10194\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46572\
        );

    \I__10193\ : Span4Mux_v
    port map (
            O => \N__46599\,
            I => \N__46569\
        );

    \I__10192\ : Span4Mux_h
    port map (
            O => \N__46596\,
            I => \N__46564\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__46593\,
            I => \N__46564\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__46588\,
            I => \N__46561\
        );

    \I__10189\ : Span4Mux_h
    port map (
            O => \N__46585\,
            I => \N__46558\
        );

    \I__10188\ : Span12Mux_v
    port map (
            O => \N__46582\,
            I => \N__46555\
        );

    \I__10187\ : Span4Mux_v
    port map (
            O => \N__46575\,
            I => \N__46552\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__46572\,
            I => \N__46541\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__46569\,
            I => \N__46541\
        );

    \I__10184\ : Span4Mux_h
    port map (
            O => \N__46564\,
            I => \N__46541\
        );

    \I__10183\ : Span4Mux_h
    port map (
            O => \N__46561\,
            I => \N__46541\
        );

    \I__10182\ : Span4Mux_h
    port map (
            O => \N__46558\,
            I => \N__46541\
        );

    \I__10181\ : Odrv12
    port map (
            O => \N__46555\,
            I => comm_buf_0_7
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__46552\,
            I => comm_buf_0_7
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__46541\,
            I => comm_buf_0_7
        );

    \I__10178\ : CascadeMux
    port map (
            O => \N__46534\,
            I => \N__46531\
        );

    \I__10177\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46527\
        );

    \I__10176\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46524\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__46527\,
            I => \N__46521\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__46524\,
            I => \N__46517\
        );

    \I__10173\ : Span4Mux_h
    port map (
            O => \N__46521\,
            I => \N__46514\
        );

    \I__10172\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46511\
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__46517\,
            I => n21964
        );

    \I__10170\ : Odrv4
    port map (
            O => \N__46514\,
            I => n21964
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__46511\,
            I => n21964
        );

    \I__10168\ : CascadeMux
    port map (
            O => \N__46504\,
            I => \N__46501\
        );

    \I__10167\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46498\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__46498\,
            I => \N__46495\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__46495\,
            I => \N__46492\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__46492\,
            I => \N__46489\
        );

    \I__10163\ : Odrv4
    port map (
            O => \N__46489\,
            I => n11379
        );

    \I__10162\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46483\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__46483\,
            I => \N__46478\
        );

    \I__10160\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46475\
        );

    \I__10159\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46471\
        );

    \I__10158\ : Span4Mux_v
    port map (
            O => \N__46478\,
            I => \N__46468\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__46475\,
            I => \N__46465\
        );

    \I__10156\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46462\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__46471\,
            I => n9
        );

    \I__10154\ : Odrv4
    port map (
            O => \N__46468\,
            I => n9
        );

    \I__10153\ : Odrv4
    port map (
            O => \N__46465\,
            I => n9
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__46462\,
            I => n9
        );

    \I__10151\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46450\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__46450\,
            I => n22059
        );

    \I__10149\ : CascadeMux
    port map (
            O => \N__46447\,
            I => \N__46444\
        );

    \I__10148\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46441\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__46441\,
            I => \N__46438\
        );

    \I__10146\ : Odrv4
    port map (
            O => \N__46438\,
            I => n26_adj_1740
        );

    \I__10145\ : CascadeMux
    port map (
            O => \N__46435\,
            I => \n18850_cascade_\
        );

    \I__10144\ : CEMux
    port map (
            O => \N__46432\,
            I => \N__46428\
        );

    \I__10143\ : CEMux
    port map (
            O => \N__46431\,
            I => \N__46423\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__46428\,
            I => \N__46420\
        );

    \I__10141\ : CEMux
    port map (
            O => \N__46427\,
            I => \N__46416\
        );

    \I__10140\ : CEMux
    port map (
            O => \N__46426\,
            I => \N__46413\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__46423\,
            I => \N__46408\
        );

    \I__10138\ : Span4Mux_h
    port map (
            O => \N__46420\,
            I => \N__46408\
        );

    \I__10137\ : CEMux
    port map (
            O => \N__46419\,
            I => \N__46405\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__46416\,
            I => \N__46399\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46396\
        );

    \I__10134\ : Span4Mux_v
    port map (
            O => \N__46408\,
            I => \N__46391\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__46405\,
            I => \N__46391\
        );

    \I__10132\ : CEMux
    port map (
            O => \N__46404\,
            I => \N__46387\
        );

    \I__10131\ : CEMux
    port map (
            O => \N__46403\,
            I => \N__46384\
        );

    \I__10130\ : CEMux
    port map (
            O => \N__46402\,
            I => \N__46381\
        );

    \I__10129\ : Span4Mux_v
    port map (
            O => \N__46399\,
            I => \N__46378\
        );

    \I__10128\ : Span12Mux_h
    port map (
            O => \N__46396\,
            I => \N__46375\
        );

    \I__10127\ : Span4Mux_h
    port map (
            O => \N__46391\,
            I => \N__46372\
        );

    \I__10126\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46369\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__46387\,
            I => n13076
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__46384\,
            I => n13076
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__46381\,
            I => n13076
        );

    \I__10122\ : Odrv4
    port map (
            O => \N__46378\,
            I => n13076
        );

    \I__10121\ : Odrv12
    port map (
            O => \N__46375\,
            I => n13076
        );

    \I__10120\ : Odrv4
    port map (
            O => \N__46372\,
            I => n13076
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__46369\,
            I => n13076
        );

    \I__10118\ : SRMux
    port map (
            O => \N__46354\,
            I => \N__46345\
        );

    \I__10117\ : SRMux
    port map (
            O => \N__46353\,
            I => \N__46342\
        );

    \I__10116\ : SRMux
    port map (
            O => \N__46352\,
            I => \N__46338\
        );

    \I__10115\ : SRMux
    port map (
            O => \N__46351\,
            I => \N__46335\
        );

    \I__10114\ : SRMux
    port map (
            O => \N__46350\,
            I => \N__46332\
        );

    \I__10113\ : SRMux
    port map (
            O => \N__46349\,
            I => \N__46329\
        );

    \I__10112\ : SRMux
    port map (
            O => \N__46348\,
            I => \N__46326\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46323\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__46342\,
            I => \N__46320\
        );

    \I__10109\ : SRMux
    port map (
            O => \N__46341\,
            I => \N__46317\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__46338\,
            I => \N__46314\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46311\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46306\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__46329\,
            I => \N__46306\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__46326\,
            I => \N__46303\
        );

    \I__10103\ : Span4Mux_h
    port map (
            O => \N__46323\,
            I => \N__46300\
        );

    \I__10102\ : Span4Mux_v
    port map (
            O => \N__46320\,
            I => \N__46297\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__46317\,
            I => \N__46290\
        );

    \I__10100\ : Span4Mux_h
    port map (
            O => \N__46314\,
            I => \N__46290\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__46311\,
            I => \N__46290\
        );

    \I__10098\ : Span4Mux_h
    port map (
            O => \N__46306\,
            I => \N__46285\
        );

    \I__10097\ : Span4Mux_h
    port map (
            O => \N__46303\,
            I => \N__46285\
        );

    \I__10096\ : Odrv4
    port map (
            O => \N__46300\,
            I => n15531
        );

    \I__10095\ : Odrv4
    port map (
            O => \N__46297\,
            I => n15531
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__46290\,
            I => n15531
        );

    \I__10093\ : Odrv4
    port map (
            O => \N__46285\,
            I => n15531
        );

    \I__10092\ : InMux
    port map (
            O => \N__46276\,
            I => \N__46273\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__46273\,
            I => \N__46270\
        );

    \I__10090\ : Span4Mux_v
    port map (
            O => \N__46270\,
            I => \N__46267\
        );

    \I__10089\ : Span4Mux_v
    port map (
            O => \N__46267\,
            I => \N__46264\
        );

    \I__10088\ : Sp12to4
    port map (
            O => \N__46264\,
            I => \N__46261\
        );

    \I__10087\ : Odrv12
    port map (
            O => \N__46261\,
            I => comm_buf_3_3
        );

    \I__10086\ : InMux
    port map (
            O => \N__46258\,
            I => \N__46254\
        );

    \I__10085\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46251\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__46254\,
            I => \N__46248\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__46251\,
            I => \N__46245\
        );

    \I__10082\ : Span4Mux_v
    port map (
            O => \N__46248\,
            I => \N__46242\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__46245\,
            I => comm_buf_6_3
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__46242\,
            I => comm_buf_6_3
        );

    \I__10079\ : InMux
    port map (
            O => \N__46237\,
            I => \N__46234\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__46234\,
            I => \N__46231\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__46231\,
            I => n18851
        );

    \I__10076\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46225\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__46225\,
            I => \N__46222\
        );

    \I__10074\ : Odrv4
    port map (
            O => \N__46222\,
            I => comm_buf_5_3
        );

    \I__10073\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46216\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__46216\,
            I => n22346
        );

    \I__10071\ : CascadeMux
    port map (
            O => \N__46213\,
            I => \n18853_cascade_\
        );

    \I__10070\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46207\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__46207\,
            I => n23378
        );

    \I__10068\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46196\
        );

    \I__10067\ : InMux
    port map (
            O => \N__46203\,
            I => \N__46192\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46189\
        );

    \I__10065\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46186\
        );

    \I__10064\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46183\
        );

    \I__10063\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46180\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46177\
        );

    \I__10061\ : InMux
    port map (
            O => \N__46195\,
            I => \N__46174\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__46192\,
            I => \N__46171\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__46189\,
            I => \N__46168\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__46186\,
            I => \N__46165\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__46183\,
            I => \N__46160\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__46180\,
            I => \N__46157\
        );

    \I__10055\ : Span4Mux_h
    port map (
            O => \N__46177\,
            I => \N__46150\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__46174\,
            I => \N__46150\
        );

    \I__10053\ : Span4Mux_h
    port map (
            O => \N__46171\,
            I => \N__46150\
        );

    \I__10052\ : Span4Mux_h
    port map (
            O => \N__46168\,
            I => \N__46145\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__46165\,
            I => \N__46145\
        );

    \I__10050\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46142\
        );

    \I__10049\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46139\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__46160\,
            I => \N__46132\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__46157\,
            I => \N__46132\
        );

    \I__10046\ : Span4Mux_v
    port map (
            O => \N__46150\,
            I => \N__46132\
        );

    \I__10045\ : Odrv4
    port map (
            O => \N__46145\,
            I => n6776
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__46142\,
            I => n6776
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__46139\,
            I => n6776
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__46132\,
            I => n6776
        );

    \I__10041\ : CascadeMux
    port map (
            O => \N__46123\,
            I => \N__46120\
        );

    \I__10040\ : InMux
    port map (
            O => \N__46120\,
            I => \N__46117\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__46117\,
            I => \N__46113\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__46116\,
            I => \N__46110\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__46113\,
            I => \N__46106\
        );

    \I__10036\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46101\
        );

    \I__10035\ : InMux
    port map (
            O => \N__46109\,
            I => \N__46101\
        );

    \I__10034\ : Sp12to4
    port map (
            O => \N__46106\,
            I => \N__46096\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__46101\,
            I => \N__46096\
        );

    \I__10032\ : Odrv12
    port map (
            O => \N__46096\,
            I => comm_buf_2_3
        );

    \I__10031\ : InMux
    port map (
            O => \N__46093\,
            I => \N__46090\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__46090\,
            I => \N__46087\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__46087\,
            I => \N__46084\
        );

    \I__10028\ : Span4Mux_h
    port map (
            O => \N__46084\,
            I => \N__46081\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__46081\,
            I => n18858
        );

    \I__10026\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46075\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__10024\ : Span4Mux_v
    port map (
            O => \N__46072\,
            I => \N__46068\
        );

    \I__10023\ : InMux
    port map (
            O => \N__46071\,
            I => \N__46065\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__46068\,
            I => \N__46062\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__46065\,
            I => \N__46059\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__46062\,
            I => \N__46053\
        );

    \I__10019\ : Span4Mux_h
    port map (
            O => \N__46059\,
            I => \N__46053\
        );

    \I__10018\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46050\
        );

    \I__10017\ : Odrv4
    port map (
            O => \N__46053\,
            I => comm_tx_buf_3
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__46050\,
            I => comm_tx_buf_3
        );

    \I__10015\ : InMux
    port map (
            O => \N__46045\,
            I => \N__46042\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__46042\,
            I => \N__46039\
        );

    \I__10013\ : Span4Mux_h
    port map (
            O => \N__46039\,
            I => \N__46036\
        );

    \I__10012\ : Sp12to4
    port map (
            O => \N__46036\,
            I => \N__46033\
        );

    \I__10011\ : Span12Mux_v
    port map (
            O => \N__46033\,
            I => \N__46030\
        );

    \I__10010\ : Span12Mux_h
    port map (
            O => \N__46030\,
            I => \N__46027\
        );

    \I__10009\ : Odrv12
    port map (
            O => \N__46027\,
            I => \THERMOSTAT\
        );

    \I__10008\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46021\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__46021\,
            I => \N__46018\
        );

    \I__10006\ : Span4Mux_h
    port map (
            O => \N__46018\,
            I => \N__46015\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__46015\,
            I => buf_control_7
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__46012\,
            I => \N__46009\
        );

    \I__10003\ : InMux
    port map (
            O => \N__46009\,
            I => \N__46002\
        );

    \I__10002\ : InMux
    port map (
            O => \N__46008\,
            I => \N__46002\
        );

    \I__10001\ : InMux
    port map (
            O => \N__46007\,
            I => \N__45999\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45992\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__45999\,
            I => \N__45989\
        );

    \I__9998\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45986\
        );

    \I__9997\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45981\
        );

    \I__9996\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45981\
        );

    \I__9995\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45978\
        );

    \I__9994\ : Span4Mux_v
    port map (
            O => \N__45992\,
            I => \N__45968\
        );

    \I__9993\ : Span4Mux_h
    port map (
            O => \N__45989\,
            I => \N__45968\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__45986\,
            I => \N__45968\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__45981\,
            I => \N__45968\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__45978\,
            I => \N__45965\
        );

    \I__9989\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45962\
        );

    \I__9988\ : Odrv4
    port map (
            O => \N__45968\,
            I => n12585
        );

    \I__9987\ : Odrv12
    port map (
            O => \N__45965\,
            I => n12585
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__45962\,
            I => n12585
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__45955\,
            I => \N__45950\
        );

    \I__9984\ : CascadeMux
    port map (
            O => \N__45954\,
            I => \N__45946\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__45953\,
            I => \N__45943\
        );

    \I__9982\ : InMux
    port map (
            O => \N__45950\,
            I => \N__45937\
        );

    \I__9981\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45934\
        );

    \I__9980\ : InMux
    port map (
            O => \N__45946\,
            I => \N__45930\
        );

    \I__9979\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45925\
        );

    \I__9978\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45925\
        );

    \I__9977\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45920\
        );

    \I__9976\ : InMux
    port map (
            O => \N__45940\,
            I => \N__45920\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__45937\,
            I => \N__45917\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__45934\,
            I => \N__45914\
        );

    \I__9973\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45911\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__45930\,
            I => \N__45904\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__45925\,
            I => \N__45904\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45904\
        );

    \I__9969\ : Span4Mux_h
    port map (
            O => \N__45917\,
            I => \N__45901\
        );

    \I__9968\ : Span4Mux_h
    port map (
            O => \N__45914\,
            I => \N__45898\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__45911\,
            I => \N__45891\
        );

    \I__9966\ : Span4Mux_v
    port map (
            O => \N__45904\,
            I => \N__45891\
        );

    \I__9965\ : Span4Mux_v
    port map (
            O => \N__45901\,
            I => \N__45891\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__45898\,
            I => n15238
        );

    \I__9963\ : Odrv4
    port map (
            O => \N__45891\,
            I => n15238
        );

    \I__9962\ : CEMux
    port map (
            O => \N__45886\,
            I => \N__45882\
        );

    \I__9961\ : InMux
    port map (
            O => \N__45885\,
            I => \N__45879\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__45882\,
            I => n12958
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__45879\,
            I => n12958
        );

    \I__9958\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45871\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__45871\,
            I => \N__45868\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__45868\,
            I => n22397
        );

    \I__9955\ : InMux
    port map (
            O => \N__45865\,
            I => \N__45862\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__45862\,
            I => n29_adj_1688
        );

    \I__9953\ : CascadeMux
    port map (
            O => \N__45859\,
            I => \n11402_cascade_\
        );

    \I__9952\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45853\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45850\
        );

    \I__9950\ : Odrv12
    port map (
            O => \N__45850\,
            I => \comm_state_3_N_500_2\
        );

    \I__9949\ : CascadeMux
    port map (
            O => \N__45847\,
            I => \n22375_cascade_\
        );

    \I__9948\ : InMux
    port map (
            O => \N__45844\,
            I => \N__45841\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__45841\,
            I => \N__45838\
        );

    \I__9946\ : Span4Mux_v
    port map (
            O => \N__45838\,
            I => \N__45835\
        );

    \I__9945\ : Span4Mux_h
    port map (
            O => \N__45835\,
            I => \N__45832\
        );

    \I__9944\ : Odrv4
    port map (
            O => \N__45832\,
            I => buf_data_iac_22
        );

    \I__9943\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45826\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__45826\,
            I => \N__45823\
        );

    \I__9941\ : Span4Mux_h
    port map (
            O => \N__45823\,
            I => \N__45820\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__45820\,
            I => n22297
        );

    \I__9939\ : InMux
    port map (
            O => \N__45817\,
            I => \N__45814\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__45814\,
            I => \N__45811\
        );

    \I__9937\ : Span4Mux_v
    port map (
            O => \N__45811\,
            I => \N__45806\
        );

    \I__9936\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45801\
        );

    \I__9935\ : InMux
    port map (
            O => \N__45809\,
            I => \N__45801\
        );

    \I__9934\ : Span4Mux_v
    port map (
            O => \N__45806\,
            I => \N__45794\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__45801\,
            I => \N__45791\
        );

    \I__9932\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45784\
        );

    \I__9931\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45774\
        );

    \I__9930\ : InMux
    port map (
            O => \N__45798\,
            I => \N__45774\
        );

    \I__9929\ : InMux
    port map (
            O => \N__45797\,
            I => \N__45774\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__45794\,
            I => \N__45769\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__45791\,
            I => \N__45769\
        );

    \I__9926\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45760\
        );

    \I__9925\ : InMux
    port map (
            O => \N__45789\,
            I => \N__45760\
        );

    \I__9924\ : InMux
    port map (
            O => \N__45788\,
            I => \N__45760\
        );

    \I__9923\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45760\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__45784\,
            I => \N__45757\
        );

    \I__9921\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45754\
        );

    \I__9920\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45749\
        );

    \I__9919\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45749\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__45774\,
            I => eis_state_1
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__45769\,
            I => eis_state_1
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__45760\,
            I => eis_state_1
        );

    \I__9915\ : Odrv4
    port map (
            O => \N__45757\,
            I => eis_state_1
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__45754\,
            I => eis_state_1
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__45749\,
            I => eis_state_1
        );

    \I__9912\ : SRMux
    port map (
            O => \N__45736\,
            I => \N__45733\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__45733\,
            I => \N__45730\
        );

    \I__9910\ : Odrv12
    port map (
            O => \N__45730\,
            I => n15517
        );

    \I__9909\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45724\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__45724\,
            I => \N__45721\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__45721\,
            I => \N__45718\
        );

    \I__9906\ : Odrv4
    port map (
            O => \N__45718\,
            I => comm_buf_3_5
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__45715\,
            I => \N__45711\
        );

    \I__9904\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45708\
        );

    \I__9903\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45705\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__45708\,
            I => comm_buf_6_5
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__45705\,
            I => comm_buf_6_5
        );

    \I__9900\ : InMux
    port map (
            O => \N__45700\,
            I => \N__45696\
        );

    \I__9899\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45692\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45689\
        );

    \I__9897\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45686\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__45692\,
            I => \N__45683\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__45689\,
            I => \N__45678\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__45686\,
            I => \N__45678\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__45683\,
            I => \N__45675\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__45678\,
            I => \N__45672\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__45675\,
            I => comm_buf_2_5
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__45672\,
            I => comm_buf_2_5
        );

    \I__9889\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45664\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__45664\,
            I => n18882
        );

    \I__9887\ : CascadeMux
    port map (
            O => \N__45661\,
            I => \n18883_cascade_\
        );

    \I__9886\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45654\
        );

    \I__9885\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45650\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__45654\,
            I => \N__45647\
        );

    \I__9883\ : InMux
    port map (
            O => \N__45653\,
            I => \N__45644\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__45650\,
            I => \N__45641\
        );

    \I__9881\ : Span4Mux_v
    port map (
            O => \N__45647\,
            I => \N__45636\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__45644\,
            I => \N__45636\
        );

    \I__9879\ : Span12Mux_v
    port map (
            O => \N__45641\,
            I => \N__45633\
        );

    \I__9878\ : Span4Mux_h
    port map (
            O => \N__45636\,
            I => \N__45630\
        );

    \I__9877\ : Odrv12
    port map (
            O => \N__45633\,
            I => comm_tx_buf_5
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__45630\,
            I => comm_tx_buf_5
        );

    \I__9875\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45622\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45619\
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__45619\,
            I => comm_buf_5_5
        );

    \I__9872\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45613\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__45613\,
            I => n22371
        );

    \I__9870\ : CascadeMux
    port map (
            O => \N__45610\,
            I => \n18885_cascade_\
        );

    \I__9869\ : InMux
    port map (
            O => \N__45607\,
            I => \N__45604\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__45604\,
            I => n23414
        );

    \I__9867\ : InMux
    port map (
            O => \N__45601\,
            I => \N__45598\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__45598\,
            I => \N__45595\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__45595\,
            I => \N__45592\
        );

    \I__9864\ : Span4Mux_h
    port map (
            O => \N__45592\,
            I => \N__45589\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__45589\,
            I => n22618
        );

    \I__9862\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45583\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__45583\,
            I => \N__45580\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__45580\,
            I => \N__45577\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__45577\,
            I => \N__45574\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__45574\,
            I => n8_adj_1755
        );

    \I__9857\ : CascadeMux
    port map (
            O => \N__45571\,
            I => \N__45566\
        );

    \I__9856\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45563\
        );

    \I__9855\ : InMux
    port map (
            O => \N__45569\,
            I => \N__45559\
        );

    \I__9854\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45553\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__45563\,
            I => \N__45550\
        );

    \I__9852\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45547\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__45559\,
            I => \N__45544\
        );

    \I__9850\ : InMux
    port map (
            O => \N__45558\,
            I => \N__45537\
        );

    \I__9849\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45537\
        );

    \I__9848\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45537\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45532\
        );

    \I__9846\ : Span4Mux_h
    port map (
            O => \N__45550\,
            I => \N__45532\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__45547\,
            I => \N__45527\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__45544\,
            I => \N__45527\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__45537\,
            I => n12976
        );

    \I__9842\ : Odrv4
    port map (
            O => \N__45532\,
            I => n12976
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__45527\,
            I => n12976
        );

    \I__9840\ : CascadeMux
    port map (
            O => \N__45520\,
            I => \n12976_cascade_\
        );

    \I__9839\ : CascadeMux
    port map (
            O => \N__45517\,
            I => \N__45514\
        );

    \I__9838\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45511\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__45511\,
            I => \N__45507\
        );

    \I__9836\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45504\
        );

    \I__9835\ : Span4Mux_v
    port map (
            O => \N__45507\,
            I => \N__45501\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__45504\,
            I => comm_buf_6_2
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__45501\,
            I => comm_buf_6_2
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__45496\,
            I => \n12_adj_1760_cascade_\
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__45493\,
            I => \n20834_cascade_\
        );

    \I__9830\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45487\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__45487\,
            I => n30_adj_1681
        );

    \I__9828\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45481\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__45481\,
            I => n33
        );

    \I__9826\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45475\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__45475\,
            I => n32
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__45472\,
            I => \n34_cascade_\
        );

    \I__9823\ : InMux
    port map (
            O => \N__45469\,
            I => \N__45466\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__45466\,
            I => n31_adj_1680
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__45463\,
            I => \n49_cascade_\
        );

    \I__9820\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45455\
        );

    \I__9819\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45451\
        );

    \I__9818\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45448\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__45455\,
            I => \N__45445\
        );

    \I__9816\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45442\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__45451\,
            I => \N__45437\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__45448\,
            I => \N__45437\
        );

    \I__9813\ : Odrv12
    port map (
            O => \N__45445\,
            I => \comm_spi.n24022\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__45442\,
            I => \comm_spi.n24022\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__45437\,
            I => \comm_spi.n24022\
        );

    \I__9810\ : CascadeMux
    port map (
            O => \N__45430\,
            I => \n8856_cascade_\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__45427\,
            I => \N__45423\
        );

    \I__9808\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45418\
        );

    \I__9807\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45415\
        );

    \I__9806\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45411\
        );

    \I__9805\ : InMux
    port map (
            O => \N__45421\,
            I => \N__45408\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__45418\,
            I => \N__45405\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__45415\,
            I => \N__45402\
        );

    \I__9802\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45397\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__45411\,
            I => \N__45394\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__45408\,
            I => \N__45391\
        );

    \I__9799\ : Span4Mux_v
    port map (
            O => \N__45405\,
            I => \N__45388\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__45402\,
            I => \N__45385\
        );

    \I__9797\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45380\
        );

    \I__9796\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45380\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__45397\,
            I => \N__45373\
        );

    \I__9794\ : Span4Mux_h
    port map (
            O => \N__45394\,
            I => \N__45373\
        );

    \I__9793\ : Span4Mux_v
    port map (
            O => \N__45391\,
            I => \N__45373\
        );

    \I__9792\ : Span4Mux_v
    port map (
            O => \N__45388\,
            I => \N__45369\
        );

    \I__9791\ : Span4Mux_v
    port map (
            O => \N__45385\,
            I => \N__45366\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__45380\,
            I => \N__45361\
        );

    \I__9789\ : Span4Mux_h
    port map (
            O => \N__45373\,
            I => \N__45361\
        );

    \I__9788\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45358\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__45369\,
            I => \N__45355\
        );

    \I__9786\ : Span4Mux_v
    port map (
            O => \N__45366\,
            I => \N__45352\
        );

    \I__9785\ : Span4Mux_v
    port map (
            O => \N__45361\,
            I => \N__45349\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__45358\,
            I => n13273
        );

    \I__9783\ : Odrv4
    port map (
            O => \N__45355\,
            I => n13273
        );

    \I__9782\ : Odrv4
    port map (
            O => \N__45352\,
            I => n13273
        );

    \I__9781\ : Odrv4
    port map (
            O => \N__45349\,
            I => n13273
        );

    \I__9780\ : CascadeMux
    port map (
            O => \N__45340\,
            I => \N__45336\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__45339\,
            I => \N__45332\
        );

    \I__9778\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45329\
        );

    \I__9777\ : InMux
    port map (
            O => \N__45335\,
            I => \N__45322\
        );

    \I__9776\ : InMux
    port map (
            O => \N__45332\,
            I => \N__45319\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__45329\,
            I => \N__45316\
        );

    \I__9774\ : CascadeMux
    port map (
            O => \N__45328\,
            I => \N__45313\
        );

    \I__9773\ : InMux
    port map (
            O => \N__45327\,
            I => \N__45309\
        );

    \I__9772\ : InMux
    port map (
            O => \N__45326\,
            I => \N__45304\
        );

    \I__9771\ : InMux
    port map (
            O => \N__45325\,
            I => \N__45304\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__45322\,
            I => \N__45301\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__45319\,
            I => \N__45298\
        );

    \I__9768\ : Span4Mux_v
    port map (
            O => \N__45316\,
            I => \N__45295\
        );

    \I__9767\ : InMux
    port map (
            O => \N__45313\,
            I => \N__45292\
        );

    \I__9766\ : InMux
    port map (
            O => \N__45312\,
            I => \N__45289\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__45309\,
            I => \N__45284\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__45304\,
            I => \N__45284\
        );

    \I__9763\ : Span4Mux_v
    port map (
            O => \N__45301\,
            I => \N__45276\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__45298\,
            I => \N__45276\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__45295\,
            I => \N__45276\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__45292\,
            I => \N__45273\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__45289\,
            I => \N__45270\
        );

    \I__9758\ : Span4Mux_v
    port map (
            O => \N__45284\,
            I => \N__45267\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45264\
        );

    \I__9756\ : Sp12to4
    port map (
            O => \N__45276\,
            I => \N__45259\
        );

    \I__9755\ : Span12Mux_v
    port map (
            O => \N__45273\,
            I => \N__45259\
        );

    \I__9754\ : Span4Mux_v
    port map (
            O => \N__45270\,
            I => \N__45254\
        );

    \I__9753\ : Span4Mux_v
    port map (
            O => \N__45267\,
            I => \N__45254\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__45264\,
            I => comm_buf_0_5
        );

    \I__9751\ : Odrv12
    port map (
            O => \N__45259\,
            I => comm_buf_0_5
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__45254\,
            I => comm_buf_0_5
        );

    \I__9749\ : CascadeMux
    port map (
            O => \N__45247\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__9748\ : InMux
    port map (
            O => \N__45244\,
            I => \N__45241\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__45241\,
            I => \comm_spi.n24019\
        );

    \I__9746\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45235\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__45235\,
            I => \comm_spi.n15344\
        );

    \I__9744\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45229\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__45229\,
            I => \comm_spi.n15345\
        );

    \I__9742\ : CascadeMux
    port map (
            O => \N__45226\,
            I => \comm_spi.n24019_cascade_\
        );

    \I__9741\ : InMux
    port map (
            O => \N__45223\,
            I => \N__45219\
        );

    \I__9740\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45216\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__45219\,
            I => \N__45211\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45216\,
            I => \N__45211\
        );

    \I__9737\ : Odrv4
    port map (
            O => \N__45211\,
            I => secclk_cnt_0
        );

    \I__9736\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45204\
        );

    \I__9735\ : InMux
    port map (
            O => \N__45207\,
            I => \N__45201\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__45204\,
            I => \N__45198\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__45201\,
            I => \N__45193\
        );

    \I__9732\ : Span4Mux_v
    port map (
            O => \N__45198\,
            I => \N__45193\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__45193\,
            I => secclk_cnt_18
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__45190\,
            I => \N__45187\
        );

    \I__9729\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45184\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45180\
        );

    \I__9727\ : InMux
    port map (
            O => \N__45183\,
            I => \N__45177\
        );

    \I__9726\ : Span4Mux_h
    port map (
            O => \N__45180\,
            I => \N__45174\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__45177\,
            I => secclk_cnt_11
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__45174\,
            I => secclk_cnt_11
        );

    \I__9723\ : InMux
    port map (
            O => \N__45169\,
            I => \N__45165\
        );

    \I__9722\ : InMux
    port map (
            O => \N__45168\,
            I => \N__45162\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__45165\,
            I => \N__45159\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__45162\,
            I => secclk_cnt_4
        );

    \I__9719\ : Odrv4
    port map (
            O => \N__45159\,
            I => secclk_cnt_4
        );

    \I__9718\ : InMux
    port map (
            O => \N__45154\,
            I => \N__45151\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__45151\,
            I => n28
        );

    \I__9716\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45144\
        );

    \I__9715\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45141\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__45144\,
            I => \N__45136\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__45141\,
            I => \N__45136\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__45136\,
            I => \N__45132\
        );

    \I__9711\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45129\
        );

    \I__9710\ : Span4Mux_v
    port map (
            O => \N__45132\,
            I => \N__45126\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__45129\,
            I => data_index_6
        );

    \I__9708\ : Odrv4
    port map (
            O => \N__45126\,
            I => data_index_6
        );

    \I__9707\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45118\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__45118\,
            I => n8_adj_1621
        );

    \I__9705\ : CascadeMux
    port map (
            O => \N__45115\,
            I => \n8_adj_1621_cascade_\
        );

    \I__9704\ : InMux
    port map (
            O => \N__45112\,
            I => \N__45106\
        );

    \I__9703\ : InMux
    port map (
            O => \N__45111\,
            I => \N__45106\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__45106\,
            I => \N__45103\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__45103\,
            I => \N__45100\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__45100\,
            I => n7_adj_1620
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__45097\,
            I => \N__45094\
        );

    \I__9698\ : CascadeBuf
    port map (
            O => \N__45094\,
            I => \N__45091\
        );

    \I__9697\ : CascadeMux
    port map (
            O => \N__45091\,
            I => \N__45088\
        );

    \I__9696\ : CascadeBuf
    port map (
            O => \N__45088\,
            I => \N__45085\
        );

    \I__9695\ : CascadeMux
    port map (
            O => \N__45085\,
            I => \N__45082\
        );

    \I__9694\ : CascadeBuf
    port map (
            O => \N__45082\,
            I => \N__45079\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__45079\,
            I => \N__45076\
        );

    \I__9692\ : CascadeBuf
    port map (
            O => \N__45076\,
            I => \N__45073\
        );

    \I__9691\ : CascadeMux
    port map (
            O => \N__45073\,
            I => \N__45070\
        );

    \I__9690\ : CascadeBuf
    port map (
            O => \N__45070\,
            I => \N__45067\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__45067\,
            I => \N__45064\
        );

    \I__9688\ : CascadeBuf
    port map (
            O => \N__45064\,
            I => \N__45061\
        );

    \I__9687\ : CascadeMux
    port map (
            O => \N__45061\,
            I => \N__45058\
        );

    \I__9686\ : CascadeBuf
    port map (
            O => \N__45058\,
            I => \N__45054\
        );

    \I__9685\ : CascadeMux
    port map (
            O => \N__45057\,
            I => \N__45051\
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__45054\,
            I => \N__45048\
        );

    \I__9683\ : CascadeBuf
    port map (
            O => \N__45051\,
            I => \N__45045\
        );

    \I__9682\ : CascadeBuf
    port map (
            O => \N__45048\,
            I => \N__45042\
        );

    \I__9681\ : CascadeMux
    port map (
            O => \N__45045\,
            I => \N__45039\
        );

    \I__9680\ : CascadeMux
    port map (
            O => \N__45042\,
            I => \N__45036\
        );

    \I__9679\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45033\
        );

    \I__9678\ : CascadeBuf
    port map (
            O => \N__45036\,
            I => \N__45030\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45027\
        );

    \I__9676\ : CascadeMux
    port map (
            O => \N__45030\,
            I => \N__45024\
        );

    \I__9675\ : Span12Mux_s10_h
    port map (
            O => \N__45027\,
            I => \N__45021\
        );

    \I__9674\ : InMux
    port map (
            O => \N__45024\,
            I => \N__45018\
        );

    \I__9673\ : Span12Mux_v
    port map (
            O => \N__45021\,
            I => \N__45015\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__45018\,
            I => \N__45012\
        );

    \I__9671\ : Odrv12
    port map (
            O => \N__45015\,
            I => \data_index_9_N_236_6\
        );

    \I__9670\ : Odrv12
    port map (
            O => \N__45012\,
            I => \data_index_9_N_236_6\
        );

    \I__9669\ : InMux
    port map (
            O => \N__45007\,
            I => \N__45003\
        );

    \I__9668\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45000\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__45003\,
            I => \N__44994\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__45000\,
            I => \N__44994\
        );

    \I__9665\ : InMux
    port map (
            O => \N__44999\,
            I => \N__44991\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__44994\,
            I => \N__44988\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__44991\,
            I => \N__44983\
        );

    \I__9662\ : Span4Mux_h
    port map (
            O => \N__44988\,
            I => \N__44983\
        );

    \I__9661\ : Odrv4
    port map (
            O => \N__44983\,
            I => data_index_7
        );

    \I__9660\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44977\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__44977\,
            I => \N__44974\
        );

    \I__9658\ : Odrv4
    port map (
            O => \N__44974\,
            I => n8_adj_1617
        );

    \I__9657\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44967\
        );

    \I__9656\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44964\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__44967\,
            I => \N__44959\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__44964\,
            I => \N__44959\
        );

    \I__9653\ : Span4Mux_v
    port map (
            O => \N__44959\,
            I => \N__44956\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__44956\,
            I => n7_adj_1616
        );

    \I__9651\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44949\
        );

    \I__9650\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44946\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44941\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__44946\,
            I => \N__44941\
        );

    \I__9647\ : Span4Mux_v
    port map (
            O => \N__44941\,
            I => \N__44937\
        );

    \I__9646\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44934\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__44937\,
            I => \N__44931\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__44934\,
            I => data_index_8
        );

    \I__9643\ : Odrv4
    port map (
            O => \N__44931\,
            I => data_index_8
        );

    \I__9642\ : InMux
    port map (
            O => \N__44926\,
            I => \N__44920\
        );

    \I__9641\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44920\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__44920\,
            I => n8_adj_1619
        );

    \I__9639\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44911\
        );

    \I__9638\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44911\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__44911\,
            I => \N__44908\
        );

    \I__9636\ : Span4Mux_v
    port map (
            O => \N__44908\,
            I => \N__44905\
        );

    \I__9635\ : Odrv4
    port map (
            O => \N__44905\,
            I => n7_adj_1618
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__44902\,
            I => \N__44899\
        );

    \I__9633\ : CascadeBuf
    port map (
            O => \N__44899\,
            I => \N__44896\
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__44896\,
            I => \N__44893\
        );

    \I__9631\ : CascadeBuf
    port map (
            O => \N__44893\,
            I => \N__44890\
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__44890\,
            I => \N__44887\
        );

    \I__9629\ : CascadeBuf
    port map (
            O => \N__44887\,
            I => \N__44884\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__44884\,
            I => \N__44881\
        );

    \I__9627\ : CascadeBuf
    port map (
            O => \N__44881\,
            I => \N__44878\
        );

    \I__9626\ : CascadeMux
    port map (
            O => \N__44878\,
            I => \N__44875\
        );

    \I__9625\ : CascadeBuf
    port map (
            O => \N__44875\,
            I => \N__44872\
        );

    \I__9624\ : CascadeMux
    port map (
            O => \N__44872\,
            I => \N__44869\
        );

    \I__9623\ : CascadeBuf
    port map (
            O => \N__44869\,
            I => \N__44866\
        );

    \I__9622\ : CascadeMux
    port map (
            O => \N__44866\,
            I => \N__44863\
        );

    \I__9621\ : CascadeBuf
    port map (
            O => \N__44863\,
            I => \N__44859\
        );

    \I__9620\ : CascadeMux
    port map (
            O => \N__44862\,
            I => \N__44856\
        );

    \I__9619\ : CascadeMux
    port map (
            O => \N__44859\,
            I => \N__44853\
        );

    \I__9618\ : CascadeBuf
    port map (
            O => \N__44856\,
            I => \N__44850\
        );

    \I__9617\ : CascadeBuf
    port map (
            O => \N__44853\,
            I => \N__44847\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__44850\,
            I => \N__44844\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__44847\,
            I => \N__44841\
        );

    \I__9614\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44838\
        );

    \I__9613\ : CascadeBuf
    port map (
            O => \N__44841\,
            I => \N__44835\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__44838\,
            I => \N__44832\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__44835\,
            I => \N__44829\
        );

    \I__9610\ : Span12Mux_h
    port map (
            O => \N__44832\,
            I => \N__44826\
        );

    \I__9609\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44823\
        );

    \I__9608\ : Span12Mux_v
    port map (
            O => \N__44826\,
            I => \N__44820\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__44823\,
            I => \N__44817\
        );

    \I__9606\ : Odrv12
    port map (
            O => \N__44820\,
            I => \data_index_9_N_236_7\
        );

    \I__9605\ : Odrv12
    port map (
            O => \N__44817\,
            I => \data_index_9_N_236_7\
        );

    \I__9604\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44809\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__44809\,
            I => \SIG_DDS.n22671\
        );

    \I__9602\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \N__44803\
        );

    \I__9601\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44800\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__44800\,
            I => \N__44797\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__44797\,
            I => \SIG_DDS.n10\
        );

    \I__9598\ : SRMux
    port map (
            O => \N__44794\,
            I => \N__44791\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__44791\,
            I => \N__44788\
        );

    \I__9596\ : Odrv12
    port map (
            O => \N__44788\,
            I => \comm_spi.imosi_N_841\
        );

    \I__9595\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44780\
        );

    \I__9594\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44777\
        );

    \I__9593\ : InMux
    port map (
            O => \N__44783\,
            I => \N__44774\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__44780\,
            I => \N__44769\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__44777\,
            I => \N__44769\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__44774\,
            I => \comm_spi.n15331\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__44769\,
            I => \comm_spi.n15331\
        );

    \I__9588\ : CascadeMux
    port map (
            O => \N__44764\,
            I => \N__44760\
        );

    \I__9587\ : CascadeMux
    port map (
            O => \N__44763\,
            I => \N__44756\
        );

    \I__9586\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44751\
        );

    \I__9585\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44751\
        );

    \I__9584\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44748\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__44751\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__44748\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__44743\,
            I => \N__44739\
        );

    \I__9580\ : InMux
    port map (
            O => \N__44742\,
            I => \N__44734\
        );

    \I__9579\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44729\
        );

    \I__9578\ : InMux
    port map (
            O => \N__44738\,
            I => \N__44729\
        );

    \I__9577\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44726\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__44734\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__44729\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__44726\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__44719\,
            I => \N__44716\
        );

    \I__9572\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44711\
        );

    \I__9571\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44708\
        );

    \I__9570\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44704\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44700\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__44708\,
            I => \N__44697\
        );

    \I__9567\ : CascadeMux
    port map (
            O => \N__44707\,
            I => \N__44694\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__44704\,
            I => \N__44690\
        );

    \I__9565\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44687\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__44700\,
            I => \N__44684\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__44697\,
            I => \N__44681\
        );

    \I__9562\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44678\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__44693\,
            I => \N__44674\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__44690\,
            I => \N__44665\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__44687\,
            I => \N__44665\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__44684\,
            I => \N__44665\
        );

    \I__9557\ : Span4Mux_h
    port map (
            O => \N__44681\,
            I => \N__44665\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__44678\,
            I => \N__44662\
        );

    \I__9555\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44657\
        );

    \I__9554\ : InMux
    port map (
            O => \N__44674\,
            I => \N__44657\
        );

    \I__9553\ : Span4Mux_v
    port map (
            O => \N__44665\,
            I => \N__44654\
        );

    \I__9552\ : Odrv12
    port map (
            O => \N__44662\,
            I => comm_buf_0_4
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__44657\,
            I => comm_buf_0_4
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__44654\,
            I => comm_buf_0_4
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__44647\,
            I => \N__44643\
        );

    \I__9548\ : CascadeMux
    port map (
            O => \N__44646\,
            I => \N__44639\
        );

    \I__9547\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44636\
        );

    \I__9546\ : InMux
    port map (
            O => \N__44642\,
            I => \N__44633\
        );

    \I__9545\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44627\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__44636\,
            I => \N__44624\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__44633\,
            I => \N__44621\
        );

    \I__9542\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44618\
        );

    \I__9541\ : CascadeMux
    port map (
            O => \N__44631\,
            I => \N__44614\
        );

    \I__9540\ : CascadeMux
    port map (
            O => \N__44630\,
            I => \N__44610\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__44627\,
            I => \N__44607\
        );

    \I__9538\ : Span4Mux_v
    port map (
            O => \N__44624\,
            I => \N__44604\
        );

    \I__9537\ : Span4Mux_v
    port map (
            O => \N__44621\,
            I => \N__44599\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__44618\,
            I => \N__44599\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__44617\,
            I => \N__44596\
        );

    \I__9534\ : InMux
    port map (
            O => \N__44614\,
            I => \N__44593\
        );

    \I__9533\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44589\
        );

    \I__9532\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44586\
        );

    \I__9531\ : Span4Mux_v
    port map (
            O => \N__44607\,
            I => \N__44583\
        );

    \I__9530\ : Span4Mux_v
    port map (
            O => \N__44604\,
            I => \N__44578\
        );

    \I__9529\ : Span4Mux_h
    port map (
            O => \N__44599\,
            I => \N__44578\
        );

    \I__9528\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44575\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__44593\,
            I => \N__44572\
        );

    \I__9526\ : InMux
    port map (
            O => \N__44592\,
            I => \N__44569\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__44589\,
            I => \N__44566\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__44586\,
            I => \N__44558\
        );

    \I__9523\ : Span4Mux_h
    port map (
            O => \N__44583\,
            I => \N__44558\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__44578\,
            I => \N__44558\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__44575\,
            I => \N__44555\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__44572\,
            I => \N__44552\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__44569\,
            I => \N__44549\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__44566\,
            I => \N__44546\
        );

    \I__9517\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44543\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__44558\,
            I => \N__44540\
        );

    \I__9515\ : Odrv12
    port map (
            O => \N__44555\,
            I => comm_buf_0_1
        );

    \I__9514\ : Odrv4
    port map (
            O => \N__44552\,
            I => comm_buf_0_1
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__44549\,
            I => comm_buf_0_1
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__44546\,
            I => comm_buf_0_1
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__44543\,
            I => comm_buf_0_1
        );

    \I__9510\ : Odrv4
    port map (
            O => \N__44540\,
            I => comm_buf_0_1
        );

    \I__9509\ : InMux
    port map (
            O => \N__44527\,
            I => \N__44523\
        );

    \I__9508\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44520\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__44523\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__44520\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__9505\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44509\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__44509\,
            I => \N__44505\
        );

    \I__9502\ : InMux
    port map (
            O => \N__44508\,
            I => \N__44502\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__44505\,
            I => n8_adj_1615
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__44502\,
            I => n8_adj_1615
        );

    \I__9499\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44493\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44490\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__44493\,
            I => \N__44487\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__44490\,
            I => \N__44484\
        );

    \I__9495\ : Span4Mux_v
    port map (
            O => \N__44487\,
            I => \N__44479\
        );

    \I__9494\ : Span4Mux_v
    port map (
            O => \N__44484\,
            I => \N__44479\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__44479\,
            I => n7_adj_1614
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__44476\,
            I => \N__44473\
        );

    \I__9491\ : CascadeBuf
    port map (
            O => \N__44473\,
            I => \N__44470\
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__44470\,
            I => \N__44467\
        );

    \I__9489\ : CascadeBuf
    port map (
            O => \N__44467\,
            I => \N__44464\
        );

    \I__9488\ : CascadeMux
    port map (
            O => \N__44464\,
            I => \N__44461\
        );

    \I__9487\ : CascadeBuf
    port map (
            O => \N__44461\,
            I => \N__44458\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__44458\,
            I => \N__44455\
        );

    \I__9485\ : CascadeBuf
    port map (
            O => \N__44455\,
            I => \N__44452\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__44452\,
            I => \N__44449\
        );

    \I__9483\ : CascadeBuf
    port map (
            O => \N__44449\,
            I => \N__44446\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__44446\,
            I => \N__44443\
        );

    \I__9481\ : CascadeBuf
    port map (
            O => \N__44443\,
            I => \N__44440\
        );

    \I__9480\ : CascadeMux
    port map (
            O => \N__44440\,
            I => \N__44437\
        );

    \I__9479\ : CascadeBuf
    port map (
            O => \N__44437\,
            I => \N__44434\
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__44434\,
            I => \N__44430\
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__44433\,
            I => \N__44427\
        );

    \I__9476\ : CascadeBuf
    port map (
            O => \N__44430\,
            I => \N__44424\
        );

    \I__9475\ : CascadeBuf
    port map (
            O => \N__44427\,
            I => \N__44421\
        );

    \I__9474\ : CascadeMux
    port map (
            O => \N__44424\,
            I => \N__44418\
        );

    \I__9473\ : CascadeMux
    port map (
            O => \N__44421\,
            I => \N__44415\
        );

    \I__9472\ : CascadeBuf
    port map (
            O => \N__44418\,
            I => \N__44412\
        );

    \I__9471\ : InMux
    port map (
            O => \N__44415\,
            I => \N__44409\
        );

    \I__9470\ : CascadeMux
    port map (
            O => \N__44412\,
            I => \N__44406\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__44409\,
            I => \N__44403\
        );

    \I__9468\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44400\
        );

    \I__9467\ : Span12Mux_h
    port map (
            O => \N__44403\,
            I => \N__44397\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__44400\,
            I => \N__44394\
        );

    \I__9465\ : Span12Mux_v
    port map (
            O => \N__44397\,
            I => \N__44391\
        );

    \I__9464\ : Span4Mux_h
    port map (
            O => \N__44394\,
            I => \N__44388\
        );

    \I__9463\ : Odrv12
    port map (
            O => \N__44391\,
            I => \data_index_9_N_236_9\
        );

    \I__9462\ : Odrv4
    port map (
            O => \N__44388\,
            I => \data_index_9_N_236_9\
        );

    \I__9461\ : InMux
    port map (
            O => \N__44383\,
            I => \N__44378\
        );

    \I__9460\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44375\
        );

    \I__9459\ : InMux
    port map (
            O => \N__44381\,
            I => \N__44372\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__44378\,
            I => req_data_cnt_15
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__44375\,
            I => req_data_cnt_15
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__44372\,
            I => req_data_cnt_15
        );

    \I__9455\ : InMux
    port map (
            O => \N__44365\,
            I => \N__44362\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__44362\,
            I => \N__44359\
        );

    \I__9453\ : Span4Mux_h
    port map (
            O => \N__44359\,
            I => \N__44356\
        );

    \I__9452\ : Span4Mux_h
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__44353\,
            I => n22314
        );

    \I__9450\ : InMux
    port map (
            O => \N__44350\,
            I => \N__44347\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__44347\,
            I => n22169
        );

    \I__9448\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44341\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__44341\,
            I => \N__44337\
        );

    \I__9446\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44333\
        );

    \I__9445\ : Span12Mux_h
    port map (
            O => \N__44337\,
            I => \N__44330\
        );

    \I__9444\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44327\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__44333\,
            I => req_data_cnt_3
        );

    \I__9442\ : Odrv12
    port map (
            O => \N__44330\,
            I => req_data_cnt_3
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__44327\,
            I => req_data_cnt_3
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__44320\,
            I => \n23312_cascade_\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__44317\,
            I => \n23315_cascade_\
        );

    \I__9438\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44311\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44308\
        );

    \I__9436\ : Sp12to4
    port map (
            O => \N__44308\,
            I => \N__44305\
        );

    \I__9435\ : Span12Mux_v
    port map (
            O => \N__44305\,
            I => \N__44302\
        );

    \I__9434\ : Odrv12
    port map (
            O => \N__44302\,
            I => n111_adj_1744
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__44299\,
            I => \n30_adj_1741_cascade_\
        );

    \I__9432\ : CascadeMux
    port map (
            O => \N__44296\,
            I => \N__44292\
        );

    \I__9431\ : CascadeMux
    port map (
            O => \N__44295\,
            I => \N__44289\
        );

    \I__9430\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44285\
        );

    \I__9429\ : InMux
    port map (
            O => \N__44289\,
            I => \N__44280\
        );

    \I__9428\ : InMux
    port map (
            O => \N__44288\,
            I => \N__44280\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44277\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__44280\,
            I => \acadc_skipCount_3\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__44277\,
            I => \acadc_skipCount_3\
        );

    \I__9424\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44269\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__44269\,
            I => \N__44266\
        );

    \I__9422\ : Span4Mux_v
    port map (
            O => \N__44266\,
            I => \N__44263\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__44263\,
            I => n19_adj_1739
        );

    \I__9420\ : CascadeMux
    port map (
            O => \N__44260\,
            I => \N__44257\
        );

    \I__9419\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44254\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__44254\,
            I => \N__44251\
        );

    \I__9417\ : Span4Mux_h
    port map (
            O => \N__44251\,
            I => \N__44248\
        );

    \I__9416\ : Sp12to4
    port map (
            O => \N__44248\,
            I => \N__44244\
        );

    \I__9415\ : CascadeMux
    port map (
            O => \N__44247\,
            I => \N__44241\
        );

    \I__9414\ : Span12Mux_v
    port map (
            O => \N__44244\,
            I => \N__44238\
        );

    \I__9413\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44235\
        );

    \I__9412\ : Odrv12
    port map (
            O => \N__44238\,
            I => \buf_readRTD_3\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__44235\,
            I => \buf_readRTD_3\
        );

    \I__9410\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44225\
        );

    \I__9409\ : InMux
    port map (
            O => \N__44229\,
            I => \N__44222\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__44228\,
            I => \N__44219\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__44225\,
            I => \N__44214\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44214\
        );

    \I__9405\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44211\
        );

    \I__9404\ : Span12Mux_h
    port map (
            O => \N__44214\,
            I => \N__44208\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__44211\,
            I => buf_adcdata_iac_11
        );

    \I__9402\ : Odrv12
    port map (
            O => \N__44208\,
            I => buf_adcdata_iac_11
        );

    \I__9401\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44200\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__44200\,
            I => \N__44197\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__44197\,
            I => \N__44194\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__44194\,
            I => n16_adj_1738
        );

    \I__9397\ : CascadeMux
    port map (
            O => \N__44191\,
            I => \n23558_cascade_\
        );

    \I__9396\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44185\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__44185\,
            I => n23561
        );

    \I__9394\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44176\
        );

    \I__9393\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44176\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__44176\,
            I => \N__44173\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__44173\,
            I => n7_adj_1624
        );

    \I__9390\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44167\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__44167\,
            I => n8_adj_1625
        );

    \I__9388\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44160\
        );

    \I__9387\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44157\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__44160\,
            I => \N__44151\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44151\
        );

    \I__9384\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44148\
        );

    \I__9383\ : Span4Mux_h
    port map (
            O => \N__44151\,
            I => \N__44145\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__44148\,
            I => data_index_4
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__44145\,
            I => data_index_4
        );

    \I__9380\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44137\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__44137\,
            I => n23546
        );

    \I__9378\ : InMux
    port map (
            O => \N__44134\,
            I => \N__44131\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__44131\,
            I => n30
        );

    \I__9376\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44125\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__44125\,
            I => \N__44122\
        );

    \I__9374\ : Span4Mux_h
    port map (
            O => \N__44122\,
            I => \N__44119\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__44119\,
            I => n17_adj_1594
        );

    \I__9372\ : InMux
    port map (
            O => \N__44116\,
            I => \N__44112\
        );

    \I__9371\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44109\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__44112\,
            I => \N__44106\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__44109\,
            I => \N__44100\
        );

    \I__9368\ : Span4Mux_h
    port map (
            O => \N__44106\,
            I => \N__44100\
        );

    \I__9367\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44097\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__44100\,
            I => \acadc_skipCount_8\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__44097\,
            I => \acadc_skipCount_8\
        );

    \I__9364\ : CascadeMux
    port map (
            O => \N__44092\,
            I => \N__44089\
        );

    \I__9363\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44086\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__44086\,
            I => \N__44083\
        );

    \I__9361\ : Odrv4
    port map (
            O => \N__44083\,
            I => n24_adj_1800
        );

    \I__9360\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44075\
        );

    \I__9359\ : CascadeMux
    port map (
            O => \N__44079\,
            I => \N__44072\
        );

    \I__9358\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44069\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44066\
        );

    \I__9356\ : InMux
    port map (
            O => \N__44072\,
            I => \N__44063\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__44069\,
            I => req_data_cnt_9
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__44066\,
            I => req_data_cnt_9
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__44063\,
            I => req_data_cnt_9
        );

    \I__9352\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44053\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__44053\,
            I => \N__44050\
        );

    \I__9350\ : Sp12to4
    port map (
            O => \N__44050\,
            I => \N__44047\
        );

    \I__9349\ : Odrv12
    port map (
            O => \N__44047\,
            I => n18_adj_1699
        );

    \I__9348\ : CEMux
    port map (
            O => \N__44044\,
            I => \N__44041\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__44041\,
            I => \N__44037\
        );

    \I__9346\ : CascadeMux
    port map (
            O => \N__44040\,
            I => \N__44034\
        );

    \I__9345\ : Span4Mux_h
    port map (
            O => \N__44037\,
            I => \N__44031\
        );

    \I__9344\ : InMux
    port map (
            O => \N__44034\,
            I => \N__44028\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__44031\,
            I => \N__44025\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__44022\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__44025\,
            I => n13257
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__44022\,
            I => n13257
        );

    \I__9339\ : InMux
    port map (
            O => \N__44017\,
            I => \N__44014\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__44014\,
            I => \N__44011\
        );

    \I__9337\ : Span4Mux_v
    port map (
            O => \N__44011\,
            I => \N__44007\
        );

    \I__9336\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44004\
        );

    \I__9335\ : Span4Mux_h
    port map (
            O => \N__44007\,
            I => \N__44001\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__44004\,
            I => acadc_skipcnt_1
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__44001\,
            I => acadc_skipcnt_1
        );

    \I__9332\ : CascadeMux
    port map (
            O => \N__43996\,
            I => \N__43993\
        );

    \I__9331\ : InMux
    port map (
            O => \N__43993\,
            I => \N__43990\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__43990\,
            I => \N__43987\
        );

    \I__9329\ : Span4Mux_v
    port map (
            O => \N__43987\,
            I => \N__43983\
        );

    \I__9328\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43980\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__43983\,
            I => \N__43977\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__43980\,
            I => acadc_skipcnt_4
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__43977\,
            I => acadc_skipcnt_4
        );

    \I__9324\ : InMux
    port map (
            O => \N__43972\,
            I => \N__43969\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__43969\,
            I => \N__43966\
        );

    \I__9322\ : Span4Mux_h
    port map (
            O => \N__43966\,
            I => \N__43963\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__43963\,
            I => n18
        );

    \I__9320\ : InMux
    port map (
            O => \N__43960\,
            I => \N__43957\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__43957\,
            I => \N__43952\
        );

    \I__9318\ : CascadeMux
    port map (
            O => \N__43956\,
            I => \N__43949\
        );

    \I__9317\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43944\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__43952\,
            I => \N__43941\
        );

    \I__9315\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43934\
        );

    \I__9314\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43934\
        );

    \I__9313\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43930\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__43944\,
            I => \N__43927\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__43941\,
            I => \N__43924\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__43940\,
            I => \N__43921\
        );

    \I__9309\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43918\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__43934\,
            I => \N__43915\
        );

    \I__9307\ : InMux
    port map (
            O => \N__43933\,
            I => \N__43911\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__43930\,
            I => \N__43908\
        );

    \I__9305\ : Span4Mux_h
    port map (
            O => \N__43927\,
            I => \N__43905\
        );

    \I__9304\ : Span4Mux_v
    port map (
            O => \N__43924\,
            I => \N__43902\
        );

    \I__9303\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43899\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__43918\,
            I => \N__43894\
        );

    \I__9301\ : Span4Mux_h
    port map (
            O => \N__43915\,
            I => \N__43894\
        );

    \I__9300\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43891\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__43911\,
            I => \N__43886\
        );

    \I__9298\ : Span12Mux_h
    port map (
            O => \N__43908\,
            I => \N__43886\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__43905\,
            I => comm_buf_0_0
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__43902\,
            I => comm_buf_0_0
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__43899\,
            I => comm_buf_0_0
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__43894\,
            I => comm_buf_0_0
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__43891\,
            I => comm_buf_0_0
        );

    \I__9292\ : Odrv12
    port map (
            O => \N__43886\,
            I => comm_buf_0_0
        );

    \I__9291\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43869\
        );

    \I__9290\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43866\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__43869\,
            I => \N__43862\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43859\
        );

    \I__9287\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43856\
        );

    \I__9286\ : Span4Mux_v
    port map (
            O => \N__43862\,
            I => \N__43853\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__43859\,
            I => \N__43848\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__43856\,
            I => \N__43848\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__43853\,
            I => n11172
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__43848\,
            I => n11172
        );

    \I__9281\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43839\
        );

    \I__9280\ : CascadeMux
    port map (
            O => \N__43842\,
            I => \N__43836\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__43839\,
            I => \N__43832\
        );

    \I__9278\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43829\
        );

    \I__9277\ : InMux
    port map (
            O => \N__43835\,
            I => \N__43825\
        );

    \I__9276\ : Span4Mux_v
    port map (
            O => \N__43832\,
            I => \N__43822\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__43829\,
            I => \N__43819\
        );

    \I__9274\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43815\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__43825\,
            I => \N__43808\
        );

    \I__9272\ : Sp12to4
    port map (
            O => \N__43822\,
            I => \N__43808\
        );

    \I__9271\ : Span12Mux_v
    port map (
            O => \N__43819\,
            I => \N__43808\
        );

    \I__9270\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43805\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__43815\,
            I => eis_start
        );

    \I__9268\ : Odrv12
    port map (
            O => \N__43808\,
            I => eis_start
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__43805\,
            I => eis_start
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__43798\,
            I => \n8_adj_1625_cascade_\
        );

    \I__9265\ : CascadeMux
    port map (
            O => \N__43795\,
            I => \N__43792\
        );

    \I__9264\ : CascadeBuf
    port map (
            O => \N__43792\,
            I => \N__43789\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__43789\,
            I => \N__43786\
        );

    \I__9262\ : CascadeBuf
    port map (
            O => \N__43786\,
            I => \N__43783\
        );

    \I__9261\ : CascadeMux
    port map (
            O => \N__43783\,
            I => \N__43780\
        );

    \I__9260\ : CascadeBuf
    port map (
            O => \N__43780\,
            I => \N__43777\
        );

    \I__9259\ : CascadeMux
    port map (
            O => \N__43777\,
            I => \N__43774\
        );

    \I__9258\ : CascadeBuf
    port map (
            O => \N__43774\,
            I => \N__43771\
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__43771\,
            I => \N__43768\
        );

    \I__9256\ : CascadeBuf
    port map (
            O => \N__43768\,
            I => \N__43765\
        );

    \I__9255\ : CascadeMux
    port map (
            O => \N__43765\,
            I => \N__43762\
        );

    \I__9254\ : CascadeBuf
    port map (
            O => \N__43762\,
            I => \N__43759\
        );

    \I__9253\ : CascadeMux
    port map (
            O => \N__43759\,
            I => \N__43755\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__43758\,
            I => \N__43752\
        );

    \I__9251\ : CascadeBuf
    port map (
            O => \N__43755\,
            I => \N__43749\
        );

    \I__9250\ : CascadeBuf
    port map (
            O => \N__43752\,
            I => \N__43746\
        );

    \I__9249\ : CascadeMux
    port map (
            O => \N__43749\,
            I => \N__43743\
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__43746\,
            I => \N__43740\
        );

    \I__9247\ : CascadeBuf
    port map (
            O => \N__43743\,
            I => \N__43737\
        );

    \I__9246\ : InMux
    port map (
            O => \N__43740\,
            I => \N__43734\
        );

    \I__9245\ : CascadeMux
    port map (
            O => \N__43737\,
            I => \N__43731\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__43734\,
            I => \N__43728\
        );

    \I__9243\ : CascadeBuf
    port map (
            O => \N__43731\,
            I => \N__43725\
        );

    \I__9242\ : Span4Mux_h
    port map (
            O => \N__43728\,
            I => \N__43722\
        );

    \I__9241\ : CascadeMux
    port map (
            O => \N__43725\,
            I => \N__43719\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__43722\,
            I => \N__43716\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43719\,
            I => \N__43713\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__43716\,
            I => \N__43710\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__43713\,
            I => \N__43707\
        );

    \I__9236\ : Sp12to4
    port map (
            O => \N__43710\,
            I => \N__43702\
        );

    \I__9235\ : Span12Mux_s11_v
    port map (
            O => \N__43707\,
            I => \N__43702\
        );

    \I__9234\ : Odrv12
    port map (
            O => \N__43702\,
            I => \data_index_9_N_236_4\
        );

    \I__9233\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43696\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__43696\,
            I => \N__43693\
        );

    \I__9231\ : Span12Mux_h
    port map (
            O => \N__43693\,
            I => \N__43690\
        );

    \I__9230\ : Odrv12
    port map (
            O => \N__43690\,
            I => n19_adj_1722
        );

    \I__9229\ : CascadeMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__9228\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43681\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__43681\,
            I => \N__43678\
        );

    \I__9226\ : Span4Mux_v
    port map (
            O => \N__43678\,
            I => \N__43675\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__43675\,
            I => \N__43672\
        );

    \I__9224\ : Sp12to4
    port map (
            O => \N__43672\,
            I => \N__43668\
        );

    \I__9223\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43665\
        );

    \I__9222\ : Odrv12
    port map (
            O => \N__43668\,
            I => \buf_readRTD_6\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__43665\,
            I => \buf_readRTD_6\
        );

    \I__9220\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43657\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__43657\,
            I => n23288
        );

    \I__9218\ : CascadeMux
    port map (
            O => \N__43654\,
            I => \n22396_cascade_\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__43651\,
            I => \N__43647\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__43650\,
            I => \N__43644\
        );

    \I__9215\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43641\
        );

    \I__9214\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43638\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__43641\,
            I => n6
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__43638\,
            I => n6
        );

    \I__9211\ : InMux
    port map (
            O => \N__43633\,
            I => \N__43629\
        );

    \I__9210\ : InMux
    port map (
            O => \N__43632\,
            I => \N__43626\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__43629\,
            I => \N__43623\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__43626\,
            I => n22061
        );

    \I__9207\ : Odrv4
    port map (
            O => \N__43623\,
            I => n22061
        );

    \I__9206\ : InMux
    port map (
            O => \N__43618\,
            I => \N__43613\
        );

    \I__9205\ : InMux
    port map (
            O => \N__43617\,
            I => \N__43606\
        );

    \I__9204\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43606\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43603\
        );

    \I__9202\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43600\
        );

    \I__9201\ : InMux
    port map (
            O => \N__43611\,
            I => \N__43597\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__43606\,
            I => \N__43592\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__43603\,
            I => \N__43592\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__43600\,
            I => \N__43589\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43586\
        );

    \I__9196\ : Span4Mux_h
    port map (
            O => \N__43592\,
            I => \N__43583\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__43589\,
            I => \N__43578\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__43586\,
            I => \N__43578\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__43583\,
            I => n21929
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__43578\,
            I => n21929
        );

    \I__9191\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43570\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__43570\,
            I => n22_adj_1801
        );

    \I__9189\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43564\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__43564\,
            I => \N__43561\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__43561\,
            I => \N__43558\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__43558\,
            I => n112_adj_1799
        );

    \I__9185\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43552\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__43552\,
            I => \N__43549\
        );

    \I__9183\ : Span4Mux_h
    port map (
            O => \N__43549\,
            I => \N__43546\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__43546\,
            I => \comm_buf_0_7_N_543_1\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43540\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43540\,
            I => \N__43537\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__43537\,
            I => \N__43533\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__43536\,
            I => \N__43530\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__43533\,
            I => \N__43527\
        );

    \I__9176\ : InMux
    port map (
            O => \N__43530\,
            I => \N__43524\
        );

    \I__9175\ : Odrv4
    port map (
            O => \N__43527\,
            I => buf_adcdata_vdc_16
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__43524\,
            I => buf_adcdata_vdc_16
        );

    \I__9173\ : CascadeMux
    port map (
            O => \N__43519\,
            I => \n23504_cascade_\
        );

    \I__9172\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43513\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__43513\,
            I => \N__43510\
        );

    \I__9170\ : Span4Mux_h
    port map (
            O => \N__43510\,
            I => \N__43506\
        );

    \I__9169\ : InMux
    port map (
            O => \N__43509\,
            I => \N__43503\
        );

    \I__9168\ : Span4Mux_h
    port map (
            O => \N__43506\,
            I => \N__43500\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__43503\,
            I => \N__43497\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__43500\,
            I => \N__43493\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__43497\,
            I => \N__43490\
        );

    \I__9164\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43487\
        );

    \I__9163\ : Span4Mux_h
    port map (
            O => \N__43493\,
            I => \N__43484\
        );

    \I__9162\ : Span4Mux_h
    port map (
            O => \N__43490\,
            I => \N__43481\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__43487\,
            I => buf_adcdata_vac_16
        );

    \I__9160\ : Odrv4
    port map (
            O => \N__43484\,
            I => buf_adcdata_vac_16
        );

    \I__9159\ : Odrv4
    port map (
            O => \N__43481\,
            I => buf_adcdata_vac_16
        );

    \I__9158\ : InMux
    port map (
            O => \N__43474\,
            I => \N__43471\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__43471\,
            I => \N__43468\
        );

    \I__9156\ : Span4Mux_v
    port map (
            O => \N__43468\,
            I => \N__43465\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__43465\,
            I => n22288
        );

    \I__9154\ : CEMux
    port map (
            O => \N__43462\,
            I => \N__43459\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__43459\,
            I => \N__43455\
        );

    \I__9152\ : InMux
    port map (
            O => \N__43458\,
            I => \N__43452\
        );

    \I__9151\ : Span4Mux_v
    port map (
            O => \N__43455\,
            I => \N__43447\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__43452\,
            I => \N__43447\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__43447\,
            I => n12838
        );

    \I__9148\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43441\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__43441\,
            I => \N__43438\
        );

    \I__9146\ : Odrv12
    port map (
            O => \N__43438\,
            I => n23306
        );

    \I__9145\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43432\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__43432\,
            I => \N__43429\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__43429\,
            I => n8_adj_1504
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__43426\,
            I => \n6_cascade_\
        );

    \I__9141\ : InMux
    port map (
            O => \N__43423\,
            I => \N__43419\
        );

    \I__9140\ : InMux
    port map (
            O => \N__43422\,
            I => \N__43416\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__43419\,
            I => \N__43412\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__43416\,
            I => \N__43409\
        );

    \I__9137\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43406\
        );

    \I__9136\ : Span4Mux_h
    port map (
            O => \N__43412\,
            I => \N__43403\
        );

    \I__9135\ : Span4Mux_v
    port map (
            O => \N__43409\,
            I => \N__43398\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43398\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__43403\,
            I => \N__43395\
        );

    \I__9132\ : Span4Mux_h
    port map (
            O => \N__43398\,
            I => \N__43392\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__43395\,
            I => n21938
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__43392\,
            I => n21938
        );

    \I__9129\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43384\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43381\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__43381\,
            I => \N__43378\
        );

    \I__9126\ : Span4Mux_h
    port map (
            O => \N__43378\,
            I => \N__43375\
        );

    \I__9125\ : Span4Mux_v
    port map (
            O => \N__43375\,
            I => \N__43372\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__43372\,
            I => buf_data_vac_3
        );

    \I__9123\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43366\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__43366\,
            I => \N__43363\
        );

    \I__9121\ : Span4Mux_v
    port map (
            O => \N__43363\,
            I => \N__43360\
        );

    \I__9120\ : Span4Mux_h
    port map (
            O => \N__43360\,
            I => \N__43357\
        );

    \I__9119\ : Odrv4
    port map (
            O => \N__43357\,
            I => buf_data_vac_2
        );

    \I__9118\ : InMux
    port map (
            O => \N__43354\,
            I => \N__43351\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__43351\,
            I => comm_buf_5_2
        );

    \I__9116\ : InMux
    port map (
            O => \N__43348\,
            I => \N__43345\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43342\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__43342\,
            I => \N__43339\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__43339\,
            I => \N__43336\
        );

    \I__9112\ : Odrv4
    port map (
            O => \N__43336\,
            I => buf_data_vac_1
        );

    \I__9111\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43330\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43327\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__43327\,
            I => \N__43324\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__43324\,
            I => comm_buf_5_1
        );

    \I__9107\ : CascadeMux
    port map (
            O => \N__43321\,
            I => \N__43318\
        );

    \I__9106\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__43312\,
            I => \N__43309\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__43309\,
            I => \N__43306\
        );

    \I__9102\ : Span4Mux_h
    port map (
            O => \N__43306\,
            I => \N__43302\
        );

    \I__9101\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43299\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__43302\,
            I => \buf_readRTD_8\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__43299\,
            I => \buf_readRTD_8\
        );

    \I__9098\ : InMux
    port map (
            O => \N__43294\,
            I => \N__43291\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__43291\,
            I => \N__43288\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__43288\,
            I => n18816
        );

    \I__9095\ : InMux
    port map (
            O => \N__43285\,
            I => \N__43281\
        );

    \I__9094\ : InMux
    port map (
            O => \N__43284\,
            I => \N__43278\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__43281\,
            I => \N__43274\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__43278\,
            I => \N__43271\
        );

    \I__9091\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43268\
        );

    \I__9090\ : Span4Mux_h
    port map (
            O => \N__43274\,
            I => \N__43265\
        );

    \I__9089\ : Span4Mux_h
    port map (
            O => \N__43271\,
            I => \N__43260\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43260\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__43265\,
            I => \N__43257\
        );

    \I__9086\ : Span4Mux_v
    port map (
            O => \N__43260\,
            I => \N__43254\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__43257\,
            I => comm_tx_buf_0
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__43254\,
            I => comm_tx_buf_0
        );

    \I__9083\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43246\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43243\
        );

    \I__9081\ : Odrv4
    port map (
            O => \N__43243\,
            I => comm_buf_3_0
        );

    \I__9080\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43237\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__43237\,
            I => n22338
        );

    \I__9078\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43231\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__43231\,
            I => n18815
        );

    \I__9076\ : CascadeMux
    port map (
            O => \N__43228\,
            I => \N__43223\
        );

    \I__9075\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43220\
        );

    \I__9074\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43217\
        );

    \I__9073\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43214\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__43220\,
            I => \N__43209\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__43217\,
            I => \N__43209\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__43214\,
            I => \N__43206\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__43209\,
            I => \N__43203\
        );

    \I__9068\ : Odrv12
    port map (
            O => \N__43206\,
            I => comm_buf_2_0
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__43203\,
            I => comm_buf_2_0
        );

    \I__9066\ : InMux
    port map (
            O => \N__43198\,
            I => \N__43195\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__9064\ : Span4Mux_h
    port map (
            O => \N__43192\,
            I => \N__43189\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__43189\,
            I => n18823
        );

    \I__9062\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43180\
        );

    \I__9060\ : Span4Mux_h
    port map (
            O => \N__43180\,
            I => \N__43177\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__43177\,
            I => \N__43174\
        );

    \I__9058\ : Odrv4
    port map (
            O => \N__43174\,
            I => buf_data_vac_0
        );

    \I__9057\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43168\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__43168\,
            I => comm_buf_5_0
        );

    \I__9055\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43162\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__43162\,
            I => \N__43159\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__43159\,
            I => \N__43156\
        );

    \I__9052\ : Span4Mux_v
    port map (
            O => \N__43156\,
            I => \N__43153\
        );

    \I__9051\ : Sp12to4
    port map (
            O => \N__43153\,
            I => \N__43150\
        );

    \I__9050\ : Odrv12
    port map (
            O => \N__43150\,
            I => buf_data_vac_7
        );

    \I__9049\ : InMux
    port map (
            O => \N__43147\,
            I => \N__43144\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__43144\,
            I => comm_buf_5_7
        );

    \I__9047\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43138\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__43138\,
            I => \N__43135\
        );

    \I__9045\ : Span4Mux_v
    port map (
            O => \N__43135\,
            I => \N__43132\
        );

    \I__9044\ : Sp12to4
    port map (
            O => \N__43132\,
            I => \N__43129\
        );

    \I__9043\ : Odrv12
    port map (
            O => \N__43129\,
            I => buf_data_vac_6
        );

    \I__9042\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43123\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__43123\,
            I => \N__43120\
        );

    \I__9040\ : Span4Mux_h
    port map (
            O => \N__43120\,
            I => \N__43117\
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__43117\,
            I => comm_buf_5_6
        );

    \I__9038\ : InMux
    port map (
            O => \N__43114\,
            I => \N__43111\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43108\
        );

    \I__9036\ : Span4Mux_v
    port map (
            O => \N__43108\,
            I => \N__43105\
        );

    \I__9035\ : Sp12to4
    port map (
            O => \N__43105\,
            I => \N__43102\
        );

    \I__9034\ : Odrv12
    port map (
            O => \N__43102\,
            I => buf_data_vac_5
        );

    \I__9033\ : InMux
    port map (
            O => \N__43099\,
            I => \N__43096\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__43096\,
            I => \N__43093\
        );

    \I__9031\ : Span4Mux_v
    port map (
            O => \N__43093\,
            I => \N__43090\
        );

    \I__9030\ : Sp12to4
    port map (
            O => \N__43090\,
            I => \N__43087\
        );

    \I__9029\ : Odrv12
    port map (
            O => \N__43087\,
            I => buf_data_vac_4
        );

    \I__9028\ : InMux
    port map (
            O => \N__43084\,
            I => \N__43081\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43081\,
            I => \N__43078\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__43078\,
            I => \N__43075\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__43075\,
            I => comm_buf_5_4
        );

    \I__9024\ : InMux
    port map (
            O => \N__43072\,
            I => \N__43068\
        );

    \I__9023\ : InMux
    port map (
            O => \N__43071\,
            I => \N__43065\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__43068\,
            I => comm_buf_6_7
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__43065\,
            I => comm_buf_6_7
        );

    \I__9020\ : InMux
    port map (
            O => \N__43060\,
            I => \N__43057\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__43057\,
            I => \N__43053\
        );

    \I__9018\ : InMux
    port map (
            O => \N__43056\,
            I => \N__43050\
        );

    \I__9017\ : Span4Mux_h
    port map (
            O => \N__43053\,
            I => \N__43047\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__43050\,
            I => comm_test_buf_24_17
        );

    \I__9015\ : Odrv4
    port map (
            O => \N__43047\,
            I => comm_test_buf_24_17
        );

    \I__9014\ : CascadeMux
    port map (
            O => \N__43042\,
            I => \N__43038\
        );

    \I__9013\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43035\
        );

    \I__9012\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43032\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43029\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__43032\,
            I => comm_buf_6_0
        );

    \I__9009\ : Odrv12
    port map (
            O => \N__43029\,
            I => comm_buf_6_0
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__43024\,
            I => \n18818_cascade_\
        );

    \I__9007\ : CascadeMux
    port map (
            O => \N__43021\,
            I => \n23372_cascade_\
        );

    \I__9006\ : InMux
    port map (
            O => \N__43018\,
            I => \N__43014\
        );

    \I__9005\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43011\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__43014\,
            I => secclk_cnt_20
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__43011\,
            I => secclk_cnt_20
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__43006\,
            I => \n20922_cascade_\
        );

    \I__9001\ : InMux
    port map (
            O => \N__43003\,
            I => \N__43000\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43000\,
            I => \N__42997\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__42997\,
            I => n14_adj_1678
        );

    \I__8998\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42990\
        );

    \I__8997\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42987\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__42990\,
            I => secclk_cnt_9
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__42987\,
            I => secclk_cnt_9
        );

    \I__8994\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42978\
        );

    \I__8993\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42975\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__42978\,
            I => \N__42972\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__42975\,
            I => secclk_cnt_17
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__42972\,
            I => secclk_cnt_17
        );

    \I__8989\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__42964\,
            I => n10_adj_1679
        );

    \I__8987\ : InMux
    port map (
            O => \N__42961\,
            I => \N__42957\
        );

    \I__8986\ : InMux
    port map (
            O => \N__42960\,
            I => \N__42954\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__42957\,
            I => secclk_cnt_6
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__42954\,
            I => secclk_cnt_6
        );

    \I__8983\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42945\
        );

    \I__8982\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42942\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__42945\,
            I => secclk_cnt_14
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__42942\,
            I => secclk_cnt_14
        );

    \I__8979\ : CascadeMux
    port map (
            O => \N__42937\,
            I => \N__42933\
        );

    \I__8978\ : InMux
    port map (
            O => \N__42936\,
            I => \N__42930\
        );

    \I__8977\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42927\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__42930\,
            I => secclk_cnt_10
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__42927\,
            I => secclk_cnt_10
        );

    \I__8974\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42918\
        );

    \I__8973\ : InMux
    port map (
            O => \N__42921\,
            I => \N__42915\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__42918\,
            I => secclk_cnt_3
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__42915\,
            I => secclk_cnt_3
        );

    \I__8970\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42907\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__42907\,
            I => n27
        );

    \I__8968\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42900\
        );

    \I__8967\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42897\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__42900\,
            I => secclk_cnt_16
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__42897\,
            I => secclk_cnt_16
        );

    \I__8964\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42888\
        );

    \I__8963\ : InMux
    port map (
            O => \N__42891\,
            I => \N__42885\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__42888\,
            I => secclk_cnt_7
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__42885\,
            I => secclk_cnt_7
        );

    \I__8960\ : CascadeMux
    port map (
            O => \N__42880\,
            I => \N__42876\
        );

    \I__8959\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42873\
        );

    \I__8958\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42870\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__42873\,
            I => secclk_cnt_13
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__42870\,
            I => secclk_cnt_13
        );

    \I__8955\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42861\
        );

    \I__8954\ : InMux
    port map (
            O => \N__42864\,
            I => \N__42858\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__42861\,
            I => secclk_cnt_2
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__42858\,
            I => secclk_cnt_2
        );

    \I__8951\ : InMux
    port map (
            O => \N__42853\,
            I => \N__42850\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__42850\,
            I => n26_adj_1715
        );

    \I__8949\ : SRMux
    port map (
            O => \N__42847\,
            I => \N__42842\
        );

    \I__8948\ : SRMux
    port map (
            O => \N__42846\,
            I => \N__42839\
        );

    \I__8947\ : SRMux
    port map (
            O => \N__42845\,
            I => \N__42836\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__42842\,
            I => \N__42833\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__42839\,
            I => \N__42830\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__42836\,
            I => \N__42827\
        );

    \I__8943\ : Span4Mux_v
    port map (
            O => \N__42833\,
            I => \N__42821\
        );

    \I__8942\ : Span4Mux_v
    port map (
            O => \N__42830\,
            I => \N__42821\
        );

    \I__8941\ : Span4Mux_h
    port map (
            O => \N__42827\,
            I => \N__42818\
        );

    \I__8940\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42815\
        );

    \I__8939\ : Odrv4
    port map (
            O => \N__42821\,
            I => n15420
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__42818\,
            I => n15420
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__42815\,
            I => n15420
        );

    \I__8936\ : IoInMux
    port map (
            O => \N__42808\,
            I => \N__42805\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__42805\,
            I => \N__42802\
        );

    \I__8934\ : Span4Mux_s2_v
    port map (
            O => \N__42802\,
            I => \N__42799\
        );

    \I__8933\ : Span4Mux_h
    port map (
            O => \N__42799\,
            I => \N__42796\
        );

    \I__8932\ : Sp12to4
    port map (
            O => \N__42796\,
            I => \N__42793\
        );

    \I__8931\ : Span12Mux_h
    port map (
            O => \N__42793\,
            I => \N__42789\
        );

    \I__8930\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42786\
        );

    \I__8929\ : Odrv12
    port map (
            O => \N__42789\,
            I => \TEST_LED\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__42786\,
            I => \TEST_LED\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__42781\,
            I => \N__42778\
        );

    \I__8926\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42775\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__42775\,
            I => \N__42772\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__42772\,
            I => \N__42769\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__42769\,
            I => n9_adj_1596
        );

    \I__8922\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42763\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__42763\,
            I => \comm_spi.n15327\
        );

    \I__8920\ : IoInMux
    port map (
            O => \N__42760\,
            I => \N__42754\
        );

    \I__8919\ : ClkMux
    port map (
            O => \N__42759\,
            I => \N__42750\
        );

    \I__8918\ : ClkMux
    port map (
            O => \N__42758\,
            I => \N__42744\
        );

    \I__8917\ : ClkMux
    port map (
            O => \N__42757\,
            I => \N__42741\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42734\
        );

    \I__8915\ : ClkMux
    port map (
            O => \N__42753\,
            I => \N__42731\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__42750\,
            I => \N__42728\
        );

    \I__8913\ : ClkMux
    port map (
            O => \N__42749\,
            I => \N__42725\
        );

    \I__8912\ : ClkMux
    port map (
            O => \N__42748\,
            I => \N__42722\
        );

    \I__8911\ : ClkMux
    port map (
            O => \N__42747\,
            I => \N__42714\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__42744\,
            I => \N__42711\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__42741\,
            I => \N__42708\
        );

    \I__8908\ : ClkMux
    port map (
            O => \N__42740\,
            I => \N__42705\
        );

    \I__8907\ : ClkMux
    port map (
            O => \N__42739\,
            I => \N__42702\
        );

    \I__8906\ : ClkMux
    port map (
            O => \N__42738\,
            I => \N__42699\
        );

    \I__8905\ : ClkMux
    port map (
            O => \N__42737\,
            I => \N__42691\
        );

    \I__8904\ : IoSpan4Mux
    port map (
            O => \N__42734\,
            I => \N__42687\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__42731\,
            I => \N__42684\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__42728\,
            I => \N__42679\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__42725\,
            I => \N__42679\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42676\
        );

    \I__8899\ : ClkMux
    port map (
            O => \N__42721\,
            I => \N__42673\
        );

    \I__8898\ : ClkMux
    port map (
            O => \N__42720\,
            I => \N__42670\
        );

    \I__8897\ : ClkMux
    port map (
            O => \N__42719\,
            I => \N__42667\
        );

    \I__8896\ : ClkMux
    port map (
            O => \N__42718\,
            I => \N__42664\
        );

    \I__8895\ : ClkMux
    port map (
            O => \N__42717\,
            I => \N__42660\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__42714\,
            I => \N__42657\
        );

    \I__8893\ : Span4Mux_v
    port map (
            O => \N__42711\,
            I => \N__42646\
        );

    \I__8892\ : Span4Mux_h
    port map (
            O => \N__42708\,
            I => \N__42646\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__42705\,
            I => \N__42646\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42646\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__42699\,
            I => \N__42646\
        );

    \I__8888\ : ClkMux
    port map (
            O => \N__42698\,
            I => \N__42643\
        );

    \I__8887\ : ClkMux
    port map (
            O => \N__42697\,
            I => \N__42640\
        );

    \I__8886\ : ClkMux
    port map (
            O => \N__42696\,
            I => \N__42637\
        );

    \I__8885\ : ClkMux
    port map (
            O => \N__42695\,
            I => \N__42634\
        );

    \I__8884\ : ClkMux
    port map (
            O => \N__42694\,
            I => \N__42631\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__42691\,
            I => \N__42628\
        );

    \I__8882\ : ClkMux
    port map (
            O => \N__42690\,
            I => \N__42625\
        );

    \I__8881\ : Sp12to4
    port map (
            O => \N__42687\,
            I => \N__42622\
        );

    \I__8880\ : Span4Mux_v
    port map (
            O => \N__42684\,
            I => \N__42617\
        );

    \I__8879\ : Span4Mux_v
    port map (
            O => \N__42679\,
            I => \N__42617\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__42676\,
            I => \N__42606\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__42673\,
            I => \N__42606\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__42670\,
            I => \N__42606\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__42667\,
            I => \N__42606\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__42664\,
            I => \N__42606\
        );

    \I__8873\ : ClkMux
    port map (
            O => \N__42663\,
            I => \N__42603\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__42660\,
            I => \N__42600\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__42657\,
            I => \N__42593\
        );

    \I__8870\ : Span4Mux_v
    port map (
            O => \N__42646\,
            I => \N__42593\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__42643\,
            I => \N__42593\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42590\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42587\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__42634\,
            I => \N__42584\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__42631\,
            I => \N__42581\
        );

    \I__8864\ : Span4Mux_h
    port map (
            O => \N__42628\,
            I => \N__42576\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__42625\,
            I => \N__42576\
        );

    \I__8862\ : Span12Mux_s6_h
    port map (
            O => \N__42622\,
            I => \N__42573\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__42617\,
            I => \N__42570\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__42606\,
            I => \N__42565\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__42603\,
            I => \N__42565\
        );

    \I__8858\ : Span4Mux_h
    port map (
            O => \N__42600\,
            I => \N__42560\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__42593\,
            I => \N__42560\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__42590\,
            I => \N__42555\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__42587\,
            I => \N__42555\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__42584\,
            I => \N__42548\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__42581\,
            I => \N__42548\
        );

    \I__8852\ : Span4Mux_v
    port map (
            O => \N__42576\,
            I => \N__42548\
        );

    \I__8851\ : Span12Mux_h
    port map (
            O => \N__42573\,
            I => \N__42543\
        );

    \I__8850\ : Sp12to4
    port map (
            O => \N__42570\,
            I => \N__42543\
        );

    \I__8849\ : Span4Mux_h
    port map (
            O => \N__42565\,
            I => \N__42540\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__42560\,
            I => \N__42537\
        );

    \I__8847\ : Span4Mux_h
    port map (
            O => \N__42555\,
            I => \N__42534\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__42548\,
            I => \N__42531\
        );

    \I__8845\ : Odrv12
    port map (
            O => \N__42543\,
            I => \VDC_CLK\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__42540\,
            I => \VDC_CLK\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__42537\,
            I => \VDC_CLK\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__42534\,
            I => \VDC_CLK\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__42531\,
            I => \VDC_CLK\
        );

    \I__8840\ : InMux
    port map (
            O => \N__42520\,
            I => \N__42517\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__42517\,
            I => \N__42514\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__42514\,
            I => n4_adj_1676
        );

    \I__8837\ : SRMux
    port map (
            O => \N__42511\,
            I => \N__42508\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__42508\,
            I => \N__42505\
        );

    \I__8835\ : Span4Mux_v
    port map (
            O => \N__42505\,
            I => \N__42502\
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__42502\,
            I => \comm_spi.DOUT_7__N_835\
        );

    \I__8833\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42495\
        );

    \I__8832\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__42495\,
            I => \N__42484\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__42492\,
            I => \N__42484\
        );

    \I__8829\ : InMux
    port map (
            O => \N__42491\,
            I => \N__42481\
        );

    \I__8828\ : InMux
    port map (
            O => \N__42490\,
            I => \N__42478\
        );

    \I__8827\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42475\
        );

    \I__8826\ : Span4Mux_v
    port map (
            O => \N__42484\,
            I => \N__42472\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__42481\,
            I => \N__42469\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__42478\,
            I => \N__42466\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__42475\,
            I => \N__42463\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__42472\,
            I => \N__42460\
        );

    \I__8821\ : Sp12to4
    port map (
            O => \N__42469\,
            I => \N__42453\
        );

    \I__8820\ : Sp12to4
    port map (
            O => \N__42466\,
            I => \N__42453\
        );

    \I__8819\ : Sp12to4
    port map (
            O => \N__42463\,
            I => \N__42453\
        );

    \I__8818\ : Sp12to4
    port map (
            O => \N__42460\,
            I => \N__42448\
        );

    \I__8817\ : Span12Mux_v
    port map (
            O => \N__42453\,
            I => \N__42448\
        );

    \I__8816\ : Span12Mux_h
    port map (
            O => \N__42448\,
            I => \N__42445\
        );

    \I__8815\ : Odrv12
    port map (
            O => \N__42445\,
            I => \ICE_SPI_SCLK\
        );

    \I__8814\ : SRMux
    port map (
            O => \N__42442\,
            I => \N__42439\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__42439\,
            I => \N__42436\
        );

    \I__8812\ : Span4Mux_h
    port map (
            O => \N__42436\,
            I => \N__42433\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__42433\,
            I => \comm_spi.iclk_N_851\
        );

    \I__8810\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42426\
        );

    \I__8809\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42423\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__42426\,
            I => secclk_cnt_15
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__42423\,
            I => secclk_cnt_15
        );

    \I__8806\ : InMux
    port map (
            O => \N__42418\,
            I => \N__42414\
        );

    \I__8805\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42411\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__42414\,
            I => secclk_cnt_8
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__42411\,
            I => secclk_cnt_8
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__42406\,
            I => \N__42402\
        );

    \I__8801\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42399\
        );

    \I__8800\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42396\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__42399\,
            I => secclk_cnt_1
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__42396\,
            I => secclk_cnt_1
        );

    \I__8797\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42387\
        );

    \I__8796\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42384\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42387\,
            I => secclk_cnt_5
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__42384\,
            I => secclk_cnt_5
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__42379\,
            I => \n25_adj_1717_cascade_\
        );

    \I__8792\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42373\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__42373\,
            I => \N__42369\
        );

    \I__8790\ : InMux
    port map (
            O => \N__42372\,
            I => \N__42366\
        );

    \I__8789\ : Span4Mux_h
    port map (
            O => \N__42369\,
            I => \N__42363\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__42366\,
            I => comm_test_buf_24_23
        );

    \I__8787\ : Odrv4
    port map (
            O => \N__42363\,
            I => comm_test_buf_24_23
        );

    \I__8786\ : InMux
    port map (
            O => \N__42358\,
            I => \N__42355\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__42355\,
            I => \N__42352\
        );

    \I__8784\ : Span4Mux_v
    port map (
            O => \N__42352\,
            I => \N__42347\
        );

    \I__8783\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42344\
        );

    \I__8782\ : InMux
    port map (
            O => \N__42350\,
            I => \N__42341\
        );

    \I__8781\ : Odrv4
    port map (
            O => \N__42347\,
            I => buf_dds0_2
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__42344\,
            I => buf_dds0_2
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__42341\,
            I => buf_dds0_2
        );

    \I__8778\ : InMux
    port map (
            O => \N__42334\,
            I => \N__42329\
        );

    \I__8777\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42326\
        );

    \I__8776\ : InMux
    port map (
            O => \N__42332\,
            I => \N__42323\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__42329\,
            I => \N__42320\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__42326\,
            I => \N__42317\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__42323\,
            I => \N__42314\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__42320\,
            I => \N__42311\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__42317\,
            I => \N__42306\
        );

    \I__8770\ : Span4Mux_v
    port map (
            O => \N__42314\,
            I => \N__42306\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__42311\,
            I => data_index_9
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__42306\,
            I => data_index_9
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__42301\,
            I => \n8_adj_1617_cascade_\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__42298\,
            I => \N__42295\
        );

    \I__8765\ : CascadeBuf
    port map (
            O => \N__42295\,
            I => \N__42292\
        );

    \I__8764\ : CascadeMux
    port map (
            O => \N__42292\,
            I => \N__42289\
        );

    \I__8763\ : CascadeBuf
    port map (
            O => \N__42289\,
            I => \N__42286\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__42286\,
            I => \N__42283\
        );

    \I__8761\ : CascadeBuf
    port map (
            O => \N__42283\,
            I => \N__42280\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__42280\,
            I => \N__42277\
        );

    \I__8759\ : CascadeBuf
    port map (
            O => \N__42277\,
            I => \N__42274\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__42274\,
            I => \N__42271\
        );

    \I__8757\ : CascadeBuf
    port map (
            O => \N__42271\,
            I => \N__42268\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__42268\,
            I => \N__42265\
        );

    \I__8755\ : CascadeBuf
    port map (
            O => \N__42265\,
            I => \N__42262\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__42262\,
            I => \N__42259\
        );

    \I__8753\ : CascadeBuf
    port map (
            O => \N__42259\,
            I => \N__42255\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__42258\,
            I => \N__42252\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__42255\,
            I => \N__42249\
        );

    \I__8750\ : CascadeBuf
    port map (
            O => \N__42252\,
            I => \N__42246\
        );

    \I__8749\ : CascadeBuf
    port map (
            O => \N__42249\,
            I => \N__42243\
        );

    \I__8748\ : CascadeMux
    port map (
            O => \N__42246\,
            I => \N__42240\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__42243\,
            I => \N__42237\
        );

    \I__8746\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42234\
        );

    \I__8745\ : CascadeBuf
    port map (
            O => \N__42237\,
            I => \N__42231\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__42234\,
            I => \N__42228\
        );

    \I__8743\ : CascadeMux
    port map (
            O => \N__42231\,
            I => \N__42225\
        );

    \I__8742\ : Span12Mux_h
    port map (
            O => \N__42228\,
            I => \N__42222\
        );

    \I__8741\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42219\
        );

    \I__8740\ : Span12Mux_v
    port map (
            O => \N__42222\,
            I => \N__42216\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__42219\,
            I => \N__42213\
        );

    \I__8738\ : Odrv12
    port map (
            O => \N__42216\,
            I => \data_index_9_N_236_8\
        );

    \I__8737\ : Odrv12
    port map (
            O => \N__42213\,
            I => \data_index_9_N_236_8\
        );

    \I__8736\ : CEMux
    port map (
            O => \N__42208\,
            I => \N__42202\
        );

    \I__8735\ : CEMux
    port map (
            O => \N__42207\,
            I => \N__42199\
        );

    \I__8734\ : CEMux
    port map (
            O => \N__42206\,
            I => \N__42196\
        );

    \I__8733\ : CEMux
    port map (
            O => \N__42205\,
            I => \N__42193\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__42202\,
            I => \N__42190\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42187\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__42196\,
            I => \N__42182\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__42193\,
            I => \N__42182\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__42190\,
            I => \N__42179\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__42187\,
            I => \N__42176\
        );

    \I__8726\ : Span4Mux_h
    port map (
            O => \N__42182\,
            I => \N__42173\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__42179\,
            I => \SIG_DDS.n13338\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__42176\,
            I => \SIG_DDS.n13338\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__42173\,
            I => \SIG_DDS.n13338\
        );

    \I__8722\ : SRMux
    port map (
            O => \N__42166\,
            I => \N__42163\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__42163\,
            I => \N__42160\
        );

    \I__8720\ : Span4Mux_h
    port map (
            O => \N__42160\,
            I => \N__42157\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__42157\,
            I => \comm_spi.iclk_N_850\
        );

    \I__8718\ : InMux
    port map (
            O => \N__42154\,
            I => \N__42149\
        );

    \I__8717\ : InMux
    port map (
            O => \N__42153\,
            I => \N__42146\
        );

    \I__8716\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42143\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__42149\,
            I => \N__42140\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__42146\,
            I => buf_dds0_1
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__42143\,
            I => buf_dds0_1
        );

    \I__8712\ : Odrv4
    port map (
            O => \N__42140\,
            I => buf_dds0_1
        );

    \I__8711\ : InMux
    port map (
            O => \N__42133\,
            I => \N__42129\
        );

    \I__8710\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42126\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__42129\,
            I => \N__42122\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__42126\,
            I => \N__42119\
        );

    \I__8707\ : InMux
    port map (
            O => \N__42125\,
            I => \N__42116\
        );

    \I__8706\ : Span4Mux_h
    port map (
            O => \N__42122\,
            I => \N__42113\
        );

    \I__8705\ : Span12Mux_s11_v
    port map (
            O => \N__42119\,
            I => \N__42110\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__42116\,
            I => buf_dds1_1
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__42113\,
            I => buf_dds1_1
        );

    \I__8702\ : Odrv12
    port map (
            O => \N__42110\,
            I => buf_dds1_1
        );

    \I__8701\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42100\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42100\,
            I => \N__42097\
        );

    \I__8699\ : Span4Mux_h
    port map (
            O => \N__42097\,
            I => \N__42092\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42089\
        );

    \I__8697\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42086\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__42092\,
            I => \N__42083\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__42089\,
            I => buf_dds1_2
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__42086\,
            I => buf_dds1_2
        );

    \I__8693\ : Odrv4
    port map (
            O => \N__42083\,
            I => buf_dds1_2
        );

    \I__8692\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42073\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__42073\,
            I => \N__42070\
        );

    \I__8690\ : Span4Mux_v
    port map (
            O => \N__42070\,
            I => \N__42066\
        );

    \I__8689\ : InMux
    port map (
            O => \N__42069\,
            I => \N__42063\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__42066\,
            I => \N__42060\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__42063\,
            I => \N__42057\
        );

    \I__8686\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42053\
        );

    \I__8685\ : Span4Mux_h
    port map (
            O => \N__42057\,
            I => \N__42050\
        );

    \I__8684\ : InMux
    port map (
            O => \N__42056\,
            I => \N__42047\
        );

    \I__8683\ : Span4Mux_h
    port map (
            O => \N__42053\,
            I => \N__42044\
        );

    \I__8682\ : Span4Mux_v
    port map (
            O => \N__42050\,
            I => \N__42041\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__42047\,
            I => buf_adcdata_iac_10
        );

    \I__8680\ : Odrv4
    port map (
            O => \N__42044\,
            I => buf_adcdata_iac_10
        );

    \I__8679\ : Odrv4
    port map (
            O => \N__42041\,
            I => buf_adcdata_iac_10
        );

    \I__8678\ : CascadeMux
    port map (
            O => \N__42034\,
            I => \n16_adj_1746_cascade_\
        );

    \I__8677\ : InMux
    port map (
            O => \N__42031\,
            I => \N__42028\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__42028\,
            I => \N__42025\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__42025\,
            I => \N__42022\
        );

    \I__8674\ : Sp12to4
    port map (
            O => \N__42022\,
            I => \N__42018\
        );

    \I__8673\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42015\
        );

    \I__8672\ : Span12Mux_v
    port map (
            O => \N__42018\,
            I => \N__42010\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__42015\,
            I => \N__42010\
        );

    \I__8670\ : Odrv12
    port map (
            O => \N__42010\,
            I => \comm_spi.n15341\
        );

    \I__8669\ : InMux
    port map (
            O => \N__42007\,
            I => \N__42004\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__42000\
        );

    \I__8667\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41997\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__42000\,
            I => \N__41994\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__41997\,
            I => \N__41991\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__41994\,
            I => \comm_spi.n15340\
        );

    \I__8663\ : Odrv12
    port map (
            O => \N__41991\,
            I => \comm_spi.n15340\
        );

    \I__8662\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41982\
        );

    \I__8661\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41977\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__41982\,
            I => \N__41974\
        );

    \I__8659\ : InMux
    port map (
            O => \N__41981\,
            I => \N__41971\
        );

    \I__8658\ : InMux
    port map (
            O => \N__41980\,
            I => \N__41967\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__41977\,
            I => \N__41964\
        );

    \I__8656\ : Span4Mux_v
    port map (
            O => \N__41974\,
            I => \N__41958\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__41971\,
            I => \N__41958\
        );

    \I__8654\ : InMux
    port map (
            O => \N__41970\,
            I => \N__41955\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__41967\,
            I => \N__41950\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__41964\,
            I => \N__41950\
        );

    \I__8651\ : InMux
    port map (
            O => \N__41963\,
            I => \N__41947\
        );

    \I__8650\ : Span4Mux_h
    port map (
            O => \N__41958\,
            I => \N__41940\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41940\
        );

    \I__8648\ : Span4Mux_v
    port map (
            O => \N__41950\,
            I => \N__41940\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__41947\,
            I => \comm_spi.n15333\
        );

    \I__8646\ : Odrv4
    port map (
            O => \N__41940\,
            I => \comm_spi.n15333\
        );

    \I__8645\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41932\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__41932\,
            I => \N__41929\
        );

    \I__8643\ : Span4Mux_v
    port map (
            O => \N__41929\,
            I => \N__41926\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__41926\,
            I => \N__41923\
        );

    \I__8641\ : Sp12to4
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__8640\ : Span12Mux_h
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__8639\ : Odrv12
    port map (
            O => \N__41917\,
            I => \comm_spi.n15334\
        );

    \I__8638\ : SRMux
    port map (
            O => \N__41914\,
            I => \N__41910\
        );

    \I__8637\ : SRMux
    port map (
            O => \N__41913\,
            I => \N__41907\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__41910\,
            I => \N__41904\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__41907\,
            I => \N__41900\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__41904\,
            I => \N__41897\
        );

    \I__8633\ : SRMux
    port map (
            O => \N__41903\,
            I => \N__41894\
        );

    \I__8632\ : Span4Mux_h
    port map (
            O => \N__41900\,
            I => \N__41891\
        );

    \I__8631\ : Span4Mux_h
    port map (
            O => \N__41897\,
            I => \N__41886\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__41894\,
            I => \N__41886\
        );

    \I__8629\ : Span4Mux_h
    port map (
            O => \N__41891\,
            I => \N__41883\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__41886\,
            I => \N__41880\
        );

    \I__8627\ : Span4Mux_v
    port map (
            O => \N__41883\,
            I => \N__41877\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__41880\,
            I => \comm_spi.data_tx_7__N_854\
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__41877\,
            I => \comm_spi.data_tx_7__N_854\
        );

    \I__8624\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41868\
        );

    \I__8623\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41864\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41861\
        );

    \I__8621\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41858\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__41864\,
            I => \N__41855\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__41861\,
            I => \N__41852\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41849\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__41855\,
            I => \N__41846\
        );

    \I__8616\ : Span4Mux_v
    port map (
            O => \N__41852\,
            I => \N__41843\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__41849\,
            I => comm_test_buf_24_1
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__41846\,
            I => comm_test_buf_24_1
        );

    \I__8613\ : Odrv4
    port map (
            O => \N__41843\,
            I => comm_test_buf_24_1
        );

    \I__8612\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41833\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__41833\,
            I => \N__41830\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__41830\,
            I => \N__41827\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__41827\,
            I => n111_adj_1798
        );

    \I__8608\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41821\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__41821\,
            I => \N__41818\
        );

    \I__8606\ : Span4Mux_v
    port map (
            O => \N__41818\,
            I => \N__41815\
        );

    \I__8605\ : Span4Mux_v
    port map (
            O => \N__41815\,
            I => \N__41812\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__41812\,
            I => n21965
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__41809\,
            I => \n12056_cascade_\
        );

    \I__8602\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41803\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__41803\,
            I => \N__41800\
        );

    \I__8600\ : Span4Mux_h
    port map (
            O => \N__41800\,
            I => \N__41797\
        );

    \I__8599\ : Span4Mux_h
    port map (
            O => \N__41797\,
            I => \N__41794\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__41794\,
            I => buf_data_iac_12
        );

    \I__8597\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41786\
        );

    \I__8596\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41783\
        );

    \I__8595\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41780\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__41786\,
            I => data_index_2
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__41783\,
            I => data_index_2
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__41780\,
            I => data_index_2
        );

    \I__8591\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41770\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__41770\,
            I => n8_adj_1628
        );

    \I__8589\ : CascadeMux
    port map (
            O => \N__41767\,
            I => \n8_adj_1628_cascade_\
        );

    \I__8588\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41758\
        );

    \I__8587\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41758\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__41758\,
            I => n7_adj_1627
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__41755\,
            I => \N__41752\
        );

    \I__8584\ : CascadeBuf
    port map (
            O => \N__41752\,
            I => \N__41749\
        );

    \I__8583\ : CascadeMux
    port map (
            O => \N__41749\,
            I => \N__41746\
        );

    \I__8582\ : CascadeBuf
    port map (
            O => \N__41746\,
            I => \N__41743\
        );

    \I__8581\ : CascadeMux
    port map (
            O => \N__41743\,
            I => \N__41740\
        );

    \I__8580\ : CascadeBuf
    port map (
            O => \N__41740\,
            I => \N__41737\
        );

    \I__8579\ : CascadeMux
    port map (
            O => \N__41737\,
            I => \N__41734\
        );

    \I__8578\ : CascadeBuf
    port map (
            O => \N__41734\,
            I => \N__41731\
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__41731\,
            I => \N__41728\
        );

    \I__8576\ : CascadeBuf
    port map (
            O => \N__41728\,
            I => \N__41725\
        );

    \I__8575\ : CascadeMux
    port map (
            O => \N__41725\,
            I => \N__41722\
        );

    \I__8574\ : CascadeBuf
    port map (
            O => \N__41722\,
            I => \N__41719\
        );

    \I__8573\ : CascadeMux
    port map (
            O => \N__41719\,
            I => \N__41715\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__41718\,
            I => \N__41712\
        );

    \I__8571\ : CascadeBuf
    port map (
            O => \N__41715\,
            I => \N__41709\
        );

    \I__8570\ : CascadeBuf
    port map (
            O => \N__41712\,
            I => \N__41706\
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__41709\,
            I => \N__41703\
        );

    \I__8568\ : CascadeMux
    port map (
            O => \N__41706\,
            I => \N__41700\
        );

    \I__8567\ : CascadeBuf
    port map (
            O => \N__41703\,
            I => \N__41697\
        );

    \I__8566\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41694\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__41697\,
            I => \N__41691\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__41694\,
            I => \N__41688\
        );

    \I__8563\ : CascadeBuf
    port map (
            O => \N__41691\,
            I => \N__41685\
        );

    \I__8562\ : Span4Mux_h
    port map (
            O => \N__41688\,
            I => \N__41682\
        );

    \I__8561\ : CascadeMux
    port map (
            O => \N__41685\,
            I => \N__41679\
        );

    \I__8560\ : Span4Mux_v
    port map (
            O => \N__41682\,
            I => \N__41676\
        );

    \I__8559\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41673\
        );

    \I__8558\ : Span4Mux_v
    port map (
            O => \N__41676\,
            I => \N__41670\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__41673\,
            I => \N__41667\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__41670\,
            I => \N__41664\
        );

    \I__8555\ : Span4Mux_h
    port map (
            O => \N__41667\,
            I => \N__41661\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__41664\,
            I => \N__41656\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__41661\,
            I => \N__41656\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__41656\,
            I => \data_index_9_N_236_2\
        );

    \I__8551\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41649\
        );

    \I__8550\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41646\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__41649\,
            I => n18865
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__41646\,
            I => n18865
        );

    \I__8547\ : InMux
    port map (
            O => \N__41641\,
            I => \N__41637\
        );

    \I__8546\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41634\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__41637\,
            I => \N__41631\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__41634\,
            I => n7_adj_1626
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__41631\,
            I => n7_adj_1626
        );

    \I__8542\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41621\
        );

    \I__8541\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41618\
        );

    \I__8540\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41615\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__41621\,
            I => data_index_3
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__41618\,
            I => data_index_3
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__41615\,
            I => data_index_3
        );

    \I__8536\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41605\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__41605\,
            I => \N__41602\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__41602\,
            I => \N__41598\
        );

    \I__8533\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41595\
        );

    \I__8532\ : Span4Mux_h
    port map (
            O => \N__41598\,
            I => \N__41592\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__41595\,
            I => acadc_skipcnt_8
        );

    \I__8530\ : Odrv4
    port map (
            O => \N__41592\,
            I => acadc_skipcnt_8
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__41587\,
            I => \N__41584\
        );

    \I__8528\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41581\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__41578\,
            I => n20
        );

    \I__8525\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41572\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__41572\,
            I => n14_adj_1599
        );

    \I__8523\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41566\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__41566\,
            I => \N__41563\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__41563\,
            I => n17
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__41560\,
            I => \n26_cascade_\
        );

    \I__8519\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41554\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__41554\,
            I => n30_adj_1743
        );

    \I__8517\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41548\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__41548\,
            I => \N__41545\
        );

    \I__8515\ : Span4Mux_h
    port map (
            O => \N__41545\,
            I => \N__41541\
        );

    \I__8514\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41538\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__41541\,
            I => n31
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__41538\,
            I => n31
        );

    \I__8511\ : InMux
    port map (
            O => \N__41533\,
            I => \N__41530\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__41530\,
            I => \N__41527\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__41527\,
            I => \N__41523\
        );

    \I__8508\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41520\
        );

    \I__8507\ : Span4Mux_v
    port map (
            O => \N__41523\,
            I => \N__41517\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__41520\,
            I => acadc_skipcnt_3
        );

    \I__8505\ : Odrv4
    port map (
            O => \N__41517\,
            I => acadc_skipcnt_3
        );

    \I__8504\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41507\
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__41511\,
            I => \N__41504\
        );

    \I__8502\ : CascadeMux
    port map (
            O => \N__41510\,
            I => \N__41501\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__41507\,
            I => \N__41498\
        );

    \I__8500\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41495\
        );

    \I__8499\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41492\
        );

    \I__8498\ : Span4Mux_h
    port map (
            O => \N__41498\,
            I => \N__41487\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__41495\,
            I => \N__41487\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__41492\,
            I => \acadc_skipCount_15\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__41487\,
            I => \acadc_skipCount_15\
        );

    \I__8494\ : InMux
    port map (
            O => \N__41482\,
            I => \N__41479\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41476\
        );

    \I__8492\ : Span4Mux_h
    port map (
            O => \N__41476\,
            I => \N__41473\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__41473\,
            I => n23_adj_1756
        );

    \I__8490\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41467\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__41467\,
            I => n21_adj_1803
        );

    \I__8488\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41461\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__41461\,
            I => \N__41458\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__41458\,
            I => n30_adj_1769
        );

    \I__8485\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41452\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__41452\,
            I => \N__41449\
        );

    \I__8483\ : Odrv4
    port map (
            O => \N__41449\,
            I => n22167
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__41446\,
            I => \N__41443\
        );

    \I__8481\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41440\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__41440\,
            I => \N__41437\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__41437\,
            I => \N__41434\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__41434\,
            I => n22166
        );

    \I__8477\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41428\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__41428\,
            I => \N__41425\
        );

    \I__8475\ : Span4Mux_h
    port map (
            O => \N__41425\,
            I => \N__41422\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__41422\,
            I => \N__41419\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__41419\,
            I => n23471
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__41416\,
            I => \n23549_cascade_\
        );

    \I__8471\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41410\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__41410\,
            I => n22174
        );

    \I__8469\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41404\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__41404\,
            I => \N__41401\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__41401\,
            I => \N__41397\
        );

    \I__8466\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41394\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__41397\,
            I => n112
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41394\,
            I => n112
        );

    \I__8463\ : InMux
    port map (
            O => \N__41389\,
            I => \N__41386\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__41386\,
            I => \N__41383\
        );

    \I__8461\ : Span4Mux_v
    port map (
            O => \N__41383\,
            I => \N__41380\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__41380\,
            I => \N__41377\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__41377\,
            I => \N__41374\
        );

    \I__8458\ : Odrv4
    port map (
            O => \N__41374\,
            I => n30_adj_1805
        );

    \I__8457\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41367\
        );

    \I__8456\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41364\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41361\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__41364\,
            I => \N__41358\
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__41361\,
            I => n17650
        );

    \I__8452\ : Odrv12
    port map (
            O => \N__41358\,
            I => n17650
        );

    \I__8451\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41350\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41346\
        );

    \I__8449\ : InMux
    port map (
            O => \N__41349\,
            I => \N__41343\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__41346\,
            I => n12
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__41343\,
            I => n12
        );

    \I__8446\ : SRMux
    port map (
            O => \N__41338\,
            I => \N__41335\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__8444\ : Span4Mux_h
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__41329\,
            I => n15553
        );

    \I__8442\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41323\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41320\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__41320\,
            I => \N__41317\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__41314\,
            I => n16_adj_1721
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__41311\,
            I => \N__41307\
        );

    \I__8436\ : InMux
    port map (
            O => \N__41310\,
            I => \N__41304\
        );

    \I__8435\ : InMux
    port map (
            O => \N__41307\,
            I => \N__41301\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__41304\,
            I => \N__41298\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__41301\,
            I => \N__41294\
        );

    \I__8432\ : Span4Mux_v
    port map (
            O => \N__41298\,
            I => \N__41291\
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__41297\,
            I => \N__41288\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__41294\,
            I => \N__41285\
        );

    \I__8429\ : Sp12to4
    port map (
            O => \N__41291\,
            I => \N__41282\
        );

    \I__8428\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41279\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__41285\,
            I => \N__41276\
        );

    \I__8426\ : Span12Mux_h
    port map (
            O => \N__41282\,
            I => \N__41273\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__41279\,
            I => buf_adcdata_iac_14
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__41276\,
            I => buf_adcdata_iac_14
        );

    \I__8423\ : Odrv12
    port map (
            O => \N__41273\,
            I => buf_adcdata_iac_14
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__41266\,
            I => \N__41262\
        );

    \I__8421\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41257\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41257\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__41257\,
            I => n12015
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__41254\,
            I => \n8_cascade_\
        );

    \I__8417\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41248\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41245\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__41245\,
            I => \N__41242\
        );

    \I__8414\ : Span4Mux_h
    port map (
            O => \N__41242\,
            I => \N__41238\
        );

    \I__8413\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41235\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__41238\,
            I => buf_adcdata_vdc_11
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__41235\,
            I => buf_adcdata_vdc_11
        );

    \I__8410\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41227\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__8408\ : Span4Mux_v
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__8407\ : Span4Mux_h
    port map (
            O => \N__41221\,
            I => \N__41217\
        );

    \I__8406\ : InMux
    port map (
            O => \N__41220\,
            I => \N__41214\
        );

    \I__8405\ : Span4Mux_h
    port map (
            O => \N__41217\,
            I => \N__41209\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41209\
        );

    \I__8403\ : Span4Mux_v
    port map (
            O => \N__41209\,
            I => \N__41205\
        );

    \I__8402\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41202\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__41205\,
            I => \N__41199\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__41202\,
            I => buf_adcdata_vac_11
        );

    \I__8399\ : Odrv4
    port map (
            O => \N__41199\,
            I => buf_adcdata_vac_11
        );

    \I__8398\ : InMux
    port map (
            O => \N__41194\,
            I => \N__41191\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__41191\,
            I => n22092
        );

    \I__8396\ : CEMux
    port map (
            O => \N__41188\,
            I => \N__41184\
        );

    \I__8395\ : InMux
    port map (
            O => \N__41187\,
            I => \N__41181\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__41184\,
            I => \N__41178\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__41181\,
            I => \N__41175\
        );

    \I__8392\ : Span12Mux_h
    port map (
            O => \N__41178\,
            I => \N__41172\
        );

    \I__8391\ : Span4Mux_h
    port map (
            O => \N__41175\,
            I => \N__41169\
        );

    \I__8390\ : Odrv12
    port map (
            O => \N__41172\,
            I => n13211
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__41169\,
            I => n13211
        );

    \I__8388\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41161\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41158\
        );

    \I__8386\ : Span4Mux_h
    port map (
            O => \N__41158\,
            I => \N__41154\
        );

    \I__8385\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41151\
        );

    \I__8384\ : Span4Mux_v
    port map (
            O => \N__41154\,
            I => \N__41148\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__41151\,
            I => acadc_skipcnt_5
        );

    \I__8382\ : Odrv4
    port map (
            O => \N__41148\,
            I => acadc_skipcnt_5
        );

    \I__8381\ : InMux
    port map (
            O => \N__41143\,
            I => \N__41140\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__41140\,
            I => \N__41137\
        );

    \I__8379\ : Span4Mux_v
    port map (
            O => \N__41137\,
            I => \N__41134\
        );

    \I__8378\ : Span4Mux_h
    port map (
            O => \N__41134\,
            I => \N__41131\
        );

    \I__8377\ : Odrv4
    port map (
            O => \N__41131\,
            I => buf_data_vac_18
        );

    \I__8376\ : InMux
    port map (
            O => \N__41128\,
            I => \N__41125\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__41125\,
            I => comm_buf_3_2
        );

    \I__8374\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41119\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__41119\,
            I => \N__41116\
        );

    \I__8372\ : Span4Mux_h
    port map (
            O => \N__41116\,
            I => \N__41113\
        );

    \I__8371\ : Span4Mux_h
    port map (
            O => \N__41113\,
            I => \N__41110\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__41110\,
            I => buf_data_vac_17
        );

    \I__8369\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41104\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__8367\ : Span4Mux_v
    port map (
            O => \N__41101\,
            I => \N__41098\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__41098\,
            I => comm_buf_3_1
        );

    \I__8365\ : SRMux
    port map (
            O => \N__41095\,
            I => \N__41092\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__41092\,
            I => \N__41089\
        );

    \I__8363\ : Span4Mux_h
    port map (
            O => \N__41089\,
            I => \N__41086\
        );

    \I__8362\ : Span4Mux_h
    port map (
            O => \N__41086\,
            I => \N__41083\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__41083\,
            I => n15503
        );

    \I__8360\ : InMux
    port map (
            O => \N__41080\,
            I => \N__41077\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__41077\,
            I => \N__41074\
        );

    \I__8358\ : Odrv12
    port map (
            O => \N__41074\,
            I => n30_adj_1708
        );

    \I__8357\ : InMux
    port map (
            O => \N__41071\,
            I => \N__41068\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__41068\,
            I => \N__41063\
        );

    \I__8355\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41058\
        );

    \I__8354\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41058\
        );

    \I__8353\ : Span12Mux_h
    port map (
            O => \N__41063\,
            I => \N__41055\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__41058\,
            I => \N__41052\
        );

    \I__8351\ : Odrv12
    port map (
            O => \N__41055\,
            I => comm_test_buf_24_2
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__41052\,
            I => comm_test_buf_24_2
        );

    \I__8349\ : InMux
    port map (
            O => \N__41047\,
            I => \N__41044\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__41044\,
            I => \N__41041\
        );

    \I__8347\ : Odrv4
    port map (
            O => \N__41041\,
            I => \comm_buf_2_7_N_575_2\
        );

    \I__8346\ : CEMux
    port map (
            O => \N__41038\,
            I => \N__41035\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__41035\,
            I => \N__41032\
        );

    \I__8344\ : Span4Mux_v
    port map (
            O => \N__41032\,
            I => \N__41028\
        );

    \I__8343\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41025\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__41028\,
            I => n12880
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__41025\,
            I => n12880
        );

    \I__8340\ : InMux
    port map (
            O => \N__41020\,
            I => \N__41016\
        );

    \I__8339\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41012\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__41016\,
            I => \N__41009\
        );

    \I__8337\ : InMux
    port map (
            O => \N__41015\,
            I => \N__41006\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__41012\,
            I => \N__41002\
        );

    \I__8335\ : Span4Mux_h
    port map (
            O => \N__41009\,
            I => \N__40997\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__41006\,
            I => \N__40997\
        );

    \I__8333\ : InMux
    port map (
            O => \N__41005\,
            I => \N__40994\
        );

    \I__8332\ : Span4Mux_h
    port map (
            O => \N__41002\,
            I => \N__40991\
        );

    \I__8331\ : Span4Mux_v
    port map (
            O => \N__40997\,
            I => \N__40986\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__40994\,
            I => \N__40986\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__40991\,
            I => n21886
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__40986\,
            I => n21886
        );

    \I__8327\ : CascadeMux
    port map (
            O => \N__40981\,
            I => \n12_cascade_\
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__40978\,
            I => \N__40975\
        );

    \I__8325\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40970\
        );

    \I__8324\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40965\
        );

    \I__8323\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40965\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__40970\,
            I => \N__40962\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__40965\,
            I => \N__40959\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__40962\,
            I => \N__40956\
        );

    \I__8319\ : Span4Mux_v
    port map (
            O => \N__40959\,
            I => \N__40953\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__40956\,
            I => comm_buf_2_2
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__40953\,
            I => comm_buf_2_2
        );

    \I__8316\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40944\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__40947\,
            I => \N__40941\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__40944\,
            I => \N__40936\
        );

    \I__8313\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40932\
        );

    \I__8312\ : InMux
    port map (
            O => \N__40940\,
            I => \N__40929\
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__40939\,
            I => \N__40926\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__40936\,
            I => \N__40921\
        );

    \I__8309\ : InMux
    port map (
            O => \N__40935\,
            I => \N__40918\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__40932\,
            I => \N__40915\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__40929\,
            I => \N__40912\
        );

    \I__8306\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40907\
        );

    \I__8305\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40907\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__40924\,
            I => \N__40904\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__40921\,
            I => \N__40899\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40899\
        );

    \I__8301\ : Span4Mux_h
    port map (
            O => \N__40915\,
            I => \N__40894\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__40912\,
            I => \N__40894\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__40907\,
            I => \N__40891\
        );

    \I__8298\ : InMux
    port map (
            O => \N__40904\,
            I => \N__40887\
        );

    \I__8297\ : Span4Mux_v
    port map (
            O => \N__40899\,
            I => \N__40884\
        );

    \I__8296\ : Span4Mux_h
    port map (
            O => \N__40894\,
            I => \N__40879\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__40891\,
            I => \N__40879\
        );

    \I__8294\ : InMux
    port map (
            O => \N__40890\,
            I => \N__40876\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__40887\,
            I => comm_buf_0_2
        );

    \I__8292\ : Odrv4
    port map (
            O => \N__40884\,
            I => comm_buf_0_2
        );

    \I__8291\ : Odrv4
    port map (
            O => \N__40879\,
            I => comm_buf_0_2
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__40876\,
            I => comm_buf_0_2
        );

    \I__8289\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40864\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__40864\,
            I => \N__40861\
        );

    \I__8287\ : Span4Mux_h
    port map (
            O => \N__40861\,
            I => \N__40858\
        );

    \I__8286\ : Odrv4
    port map (
            O => \N__40858\,
            I => n13207
        );

    \I__8285\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40849\
        );

    \I__8284\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40849\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__40849\,
            I => \N__40846\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__40846\,
            I => \N__40842\
        );

    \I__8281\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40839\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__40842\,
            I => comm_tx_buf_2
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__40839\,
            I => comm_tx_buf_2
        );

    \I__8278\ : SRMux
    port map (
            O => \N__40834\,
            I => \N__40831\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40828\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__40828\,
            I => \N__40825\
        );

    \I__8275\ : Span4Mux_v
    port map (
            O => \N__40825\,
            I => \N__40822\
        );

    \I__8274\ : Sp12to4
    port map (
            O => \N__40822\,
            I => \N__40819\
        );

    \I__8273\ : Odrv12
    port map (
            O => \N__40819\,
            I => \comm_spi.data_tx_7__N_877\
        );

    \I__8272\ : InMux
    port map (
            O => \N__40816\,
            I => \N__40813\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__8270\ : Span4Mux_h
    port map (
            O => \N__40810\,
            I => \N__40807\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__40807\,
            I => \N__40804\
        );

    \I__8268\ : Odrv4
    port map (
            O => \N__40804\,
            I => buf_data_vac_16
        );

    \I__8267\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40798\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__40798\,
            I => \N__40795\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__40795\,
            I => \N__40792\
        );

    \I__8264\ : Sp12to4
    port map (
            O => \N__40792\,
            I => \N__40789\
        );

    \I__8263\ : Span12Mux_h
    port map (
            O => \N__40789\,
            I => \N__40786\
        );

    \I__8262\ : Odrv12
    port map (
            O => \N__40786\,
            I => buf_data_vac_23
        );

    \I__8261\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40780\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__40780\,
            I => \N__40777\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__40777\,
            I => comm_buf_3_7
        );

    \I__8258\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40771\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__40771\,
            I => \N__40768\
        );

    \I__8256\ : Span4Mux_v
    port map (
            O => \N__40768\,
            I => \N__40765\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__40765\,
            I => \N__40762\
        );

    \I__8254\ : Span4Mux_h
    port map (
            O => \N__40762\,
            I => \N__40759\
        );

    \I__8253\ : Span4Mux_v
    port map (
            O => \N__40759\,
            I => \N__40756\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__40756\,
            I => buf_data_vac_22
        );

    \I__8251\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40750\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40747\
        );

    \I__8249\ : Span4Mux_v
    port map (
            O => \N__40747\,
            I => \N__40744\
        );

    \I__8248\ : Span4Mux_h
    port map (
            O => \N__40744\,
            I => \N__40741\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__40741\,
            I => comm_buf_3_6
        );

    \I__8246\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40735\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__40735\,
            I => \N__40732\
        );

    \I__8244\ : Span4Mux_h
    port map (
            O => \N__40732\,
            I => \N__40729\
        );

    \I__8243\ : Span4Mux_h
    port map (
            O => \N__40729\,
            I => \N__40726\
        );

    \I__8242\ : Span4Mux_v
    port map (
            O => \N__40726\,
            I => \N__40723\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__40723\,
            I => \N__40720\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__40720\,
            I => buf_data_vac_21
        );

    \I__8239\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40714\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__40714\,
            I => \N__40711\
        );

    \I__8237\ : Span4Mux_h
    port map (
            O => \N__40711\,
            I => \N__40708\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__40708\,
            I => \N__40705\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__40702\,
            I => buf_data_vac_20
        );

    \I__8233\ : InMux
    port map (
            O => \N__40699\,
            I => \N__40696\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__40693\,
            I => \N__40690\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__40690\,
            I => comm_buf_3_4
        );

    \I__8229\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40684\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__40684\,
            I => \N__40681\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__40681\,
            I => \N__40678\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__40678\,
            I => \N__40675\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__40675\,
            I => \N__40672\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__40672\,
            I => buf_data_vac_19
        );

    \I__8223\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40666\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__40666\,
            I => n4_adj_1664
        );

    \I__8221\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40660\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__40660\,
            I => n1
        );

    \I__8219\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40654\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__40651\,
            I => \N__40647\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__40650\,
            I => \N__40644\
        );

    \I__8215\ : Span4Mux_h
    port map (
            O => \N__40647\,
            I => \N__40640\
        );

    \I__8214\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40635\
        );

    \I__8213\ : InMux
    port map (
            O => \N__40643\,
            I => \N__40635\
        );

    \I__8212\ : Odrv4
    port map (
            O => \N__40640\,
            I => comm_tx_buf_7
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__40635\,
            I => comm_tx_buf_7
        );

    \I__8210\ : SRMux
    port map (
            O => \N__40630\,
            I => \N__40626\
        );

    \I__8209\ : SRMux
    port map (
            O => \N__40629\,
            I => \N__40623\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__40626\,
            I => \N__40620\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__40623\,
            I => \N__40616\
        );

    \I__8206\ : Span4Mux_v
    port map (
            O => \N__40620\,
            I => \N__40613\
        );

    \I__8205\ : SRMux
    port map (
            O => \N__40619\,
            I => \N__40610\
        );

    \I__8204\ : Span4Mux_v
    port map (
            O => \N__40616\,
            I => \N__40603\
        );

    \I__8203\ : Span4Mux_h
    port map (
            O => \N__40613\,
            I => \N__40603\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__40610\,
            I => \N__40603\
        );

    \I__8201\ : Span4Mux_h
    port map (
            O => \N__40603\,
            I => \N__40600\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__40600\,
            I => \comm_spi.data_tx_7__N_862\
        );

    \I__8199\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40594\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__40594\,
            I => n4_adj_1673
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__40591\,
            I => \n22342_cascade_\
        );

    \I__8196\ : InMux
    port map (
            O => \N__40588\,
            I => \N__40585\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__40585\,
            I => n23396
        );

    \I__8194\ : CascadeMux
    port map (
            O => \N__40582\,
            I => \n1_adj_1671_cascade_\
        );

    \I__8193\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8191\ : Odrv12
    port map (
            O => \N__40573\,
            I => n2_adj_1672
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__40570\,
            I => \N__40565\
        );

    \I__8189\ : CascadeMux
    port map (
            O => \N__40569\,
            I => \N__40558\
        );

    \I__8188\ : CascadeMux
    port map (
            O => \N__40568\,
            I => \N__40555\
        );

    \I__8187\ : InMux
    port map (
            O => \N__40565\,
            I => \N__40552\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__40564\,
            I => \N__40549\
        );

    \I__8185\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40546\
        );

    \I__8184\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40543\
        );

    \I__8183\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40540\
        );

    \I__8182\ : InMux
    port map (
            O => \N__40558\,
            I => \N__40536\
        );

    \I__8181\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40533\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40530\
        );

    \I__8179\ : InMux
    port map (
            O => \N__40549\,
            I => \N__40527\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__40546\,
            I => \N__40523\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__40543\,
            I => \N__40518\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40518\
        );

    \I__8175\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40514\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__40536\,
            I => \N__40509\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__40533\,
            I => \N__40509\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__40530\,
            I => \N__40504\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__40527\,
            I => \N__40504\
        );

    \I__8170\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40500\
        );

    \I__8169\ : Sp12to4
    port map (
            O => \N__40523\,
            I => \N__40497\
        );

    \I__8168\ : Span4Mux_h
    port map (
            O => \N__40518\,
            I => \N__40494\
        );

    \I__8167\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40491\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__40514\,
            I => \N__40484\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__40509\,
            I => \N__40484\
        );

    \I__8164\ : Span4Mux_h
    port map (
            O => \N__40504\,
            I => \N__40484\
        );

    \I__8163\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40481\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__40500\,
            I => \N__40476\
        );

    \I__8161\ : Span12Mux_v
    port map (
            O => \N__40497\,
            I => \N__40476\
        );

    \I__8160\ : Odrv4
    port map (
            O => \N__40494\,
            I => comm_buf_0_6
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__40491\,
            I => comm_buf_0_6
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__40484\,
            I => comm_buf_0_6
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__40481\,
            I => comm_buf_0_6
        );

    \I__8156\ : Odrv12
    port map (
            O => \N__40476\,
            I => comm_buf_0_6
        );

    \I__8155\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40462\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__40462\,
            I => \N__40458\
        );

    \I__8153\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40455\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__40458\,
            I => comm_buf_6_1
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__40455\,
            I => comm_buf_6_1
        );

    \I__8150\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40447\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__40447\,
            I => \N__40444\
        );

    \I__8148\ : Span12Mux_h
    port map (
            O => \N__40444\,
            I => \N__40441\
        );

    \I__8147\ : Odrv12
    port map (
            O => \N__40441\,
            I => buf_data_iac_2
        );

    \I__8146\ : InMux
    port map (
            O => \N__40438\,
            I => \N__40435\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__40435\,
            I => \N__40432\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__40432\,
            I => n22_adj_1707
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__40429\,
            I => \N__40426\
        );

    \I__8142\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40419\
        );

    \I__8141\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40419\
        );

    \I__8140\ : InMux
    port map (
            O => \N__40424\,
            I => \N__40416\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__40419\,
            I => \N__40413\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40410\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__40413\,
            I => \N__40407\
        );

    \I__8136\ : Span4Mux_h
    port map (
            O => \N__40410\,
            I => \N__40404\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__40407\,
            I => comm_buf_2_7
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__40404\,
            I => comm_buf_2_7
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__40399\,
            I => \n22331_cascade_\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__40396\,
            I => \n23360_cascade_\
        );

    \I__8131\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40390\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__40390\,
            I => n2_adj_1663
        );

    \I__8129\ : InMux
    port map (
            O => \N__40387\,
            I => n20806
        );

    \I__8128\ : InMux
    port map (
            O => \N__40384\,
            I => n20807
        );

    \I__8127\ : InMux
    port map (
            O => \N__40381\,
            I => n20808
        );

    \I__8126\ : InMux
    port map (
            O => \N__40378\,
            I => n20809
        );

    \I__8125\ : InMux
    port map (
            O => \N__40375\,
            I => n20810
        );

    \I__8124\ : InMux
    port map (
            O => \N__40372\,
            I => n20811
        );

    \I__8123\ : InMux
    port map (
            O => \N__40369\,
            I => \N__40365\
        );

    \I__8122\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40362\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__40365\,
            I => secclk_cnt_19
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__40362\,
            I => secclk_cnt_19
        );

    \I__8119\ : InMux
    port map (
            O => \N__40357\,
            I => \N__40353\
        );

    \I__8118\ : InMux
    port map (
            O => \N__40356\,
            I => \N__40350\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__40353\,
            I => secclk_cnt_21
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__40350\,
            I => secclk_cnt_21
        );

    \I__8115\ : CascadeMux
    port map (
            O => \N__40345\,
            I => \N__40342\
        );

    \I__8114\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40338\
        );

    \I__8113\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40335\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__40338\,
            I => \N__40332\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__40335\,
            I => secclk_cnt_12
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__40332\,
            I => secclk_cnt_12
        );

    \I__8109\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40323\
        );

    \I__8108\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40320\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__40323\,
            I => secclk_cnt_22
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__40320\,
            I => secclk_cnt_22
        );

    \I__8105\ : InMux
    port map (
            O => \N__40315\,
            I => \bfn_14_6_0_\
        );

    \I__8104\ : InMux
    port map (
            O => \N__40312\,
            I => n20798
        );

    \I__8103\ : InMux
    port map (
            O => \N__40309\,
            I => n20799
        );

    \I__8102\ : InMux
    port map (
            O => \N__40306\,
            I => n20800
        );

    \I__8101\ : InMux
    port map (
            O => \N__40303\,
            I => n20801
        );

    \I__8100\ : InMux
    port map (
            O => \N__40300\,
            I => n20802
        );

    \I__8099\ : InMux
    port map (
            O => \N__40297\,
            I => n20803
        );

    \I__8098\ : InMux
    port map (
            O => \N__40294\,
            I => n20804
        );

    \I__8097\ : InMux
    port map (
            O => \N__40291\,
            I => \bfn_14_7_0_\
        );

    \I__8096\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40284\
        );

    \I__8095\ : InMux
    port map (
            O => \N__40287\,
            I => \N__40281\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__40284\,
            I => \comm_spi.n15322\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__40281\,
            I => \comm_spi.n15322\
        );

    \I__8092\ : SRMux
    port map (
            O => \N__40276\,
            I => \N__40273\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__40273\,
            I => \N__40270\
        );

    \I__8090\ : Span4Mux_h
    port map (
            O => \N__40270\,
            I => \N__40267\
        );

    \I__8089\ : Odrv4
    port map (
            O => \N__40267\,
            I => \comm_spi.data_tx_7__N_861\
        );

    \I__8088\ : InMux
    port map (
            O => \N__40264\,
            I => \bfn_14_5_0_\
        );

    \I__8087\ : InMux
    port map (
            O => \N__40261\,
            I => n20790
        );

    \I__8086\ : InMux
    port map (
            O => \N__40258\,
            I => n20791
        );

    \I__8085\ : InMux
    port map (
            O => \N__40255\,
            I => n20792
        );

    \I__8084\ : InMux
    port map (
            O => \N__40252\,
            I => n20793
        );

    \I__8083\ : InMux
    port map (
            O => \N__40249\,
            I => n20794
        );

    \I__8082\ : InMux
    port map (
            O => \N__40246\,
            I => n20795
        );

    \I__8081\ : InMux
    port map (
            O => \N__40243\,
            I => n20796
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__40240\,
            I => \N__40237\
        );

    \I__8079\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40233\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__40236\,
            I => \N__40230\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__40233\,
            I => \N__40227\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40223\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__40227\,
            I => \N__40220\
        );

    \I__8074\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40217\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__40223\,
            I => \N__40214\
        );

    \I__8072\ : Span4Mux_v
    port map (
            O => \N__40220\,
            I => \N__40211\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__40217\,
            I => buf_dds0_8
        );

    \I__8070\ : Odrv4
    port map (
            O => \N__40214\,
            I => buf_dds0_8
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__40211\,
            I => buf_dds0_8
        );

    \I__8068\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40200\
        );

    \I__8067\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40197\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__40200\,
            I => \N__40191\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__40197\,
            I => \N__40191\
        );

    \I__8064\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40188\
        );

    \I__8063\ : Span4Mux_h
    port map (
            O => \N__40191\,
            I => \N__40185\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__40188\,
            I => data_index_1
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__40185\,
            I => data_index_1
        );

    \I__8060\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40177\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__40177\,
            I => n8_adj_1630
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \n8_adj_1630_cascade_\
        );

    \I__8057\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40165\
        );

    \I__8056\ : InMux
    port map (
            O => \N__40170\,
            I => \N__40165\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__40165\,
            I => \N__40162\
        );

    \I__8054\ : Odrv12
    port map (
            O => \N__40162\,
            I => n7_adj_1629
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__40159\,
            I => \N__40156\
        );

    \I__8052\ : CascadeBuf
    port map (
            O => \N__40156\,
            I => \N__40153\
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__40153\,
            I => \N__40150\
        );

    \I__8050\ : CascadeBuf
    port map (
            O => \N__40150\,
            I => \N__40147\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__40147\,
            I => \N__40144\
        );

    \I__8048\ : CascadeBuf
    port map (
            O => \N__40144\,
            I => \N__40141\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__40141\,
            I => \N__40138\
        );

    \I__8046\ : CascadeBuf
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__8044\ : CascadeBuf
    port map (
            O => \N__40132\,
            I => \N__40129\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__40129\,
            I => \N__40126\
        );

    \I__8042\ : CascadeBuf
    port map (
            O => \N__40126\,
            I => \N__40123\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__40123\,
            I => \N__40120\
        );

    \I__8040\ : CascadeBuf
    port map (
            O => \N__40120\,
            I => \N__40116\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__40119\,
            I => \N__40113\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__40116\,
            I => \N__40110\
        );

    \I__8037\ : CascadeBuf
    port map (
            O => \N__40113\,
            I => \N__40107\
        );

    \I__8036\ : CascadeBuf
    port map (
            O => \N__40110\,
            I => \N__40104\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \N__40101\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__40104\,
            I => \N__40098\
        );

    \I__8033\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40095\
        );

    \I__8032\ : CascadeBuf
    port map (
            O => \N__40098\,
            I => \N__40092\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__40095\,
            I => \N__40089\
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__40092\,
            I => \N__40086\
        );

    \I__8029\ : Sp12to4
    port map (
            O => \N__40089\,
            I => \N__40083\
        );

    \I__8028\ : InMux
    port map (
            O => \N__40086\,
            I => \N__40080\
        );

    \I__8027\ : Span12Mux_v
    port map (
            O => \N__40083\,
            I => \N__40077\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__40080\,
            I => \N__40074\
        );

    \I__8025\ : Odrv12
    port map (
            O => \N__40077\,
            I => \data_index_9_N_236_1\
        );

    \I__8024\ : Odrv12
    port map (
            O => \N__40074\,
            I => \data_index_9_N_236_1\
        );

    \I__8023\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40066\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__40061\
        );

    \I__8021\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40058\
        );

    \I__8020\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40055\
        );

    \I__8019\ : Span4Mux_v
    port map (
            O => \N__40061\,
            I => \N__40052\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__40058\,
            I => buf_dds0_3
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__40055\,
            I => buf_dds0_3
        );

    \I__8016\ : Odrv4
    port map (
            O => \N__40052\,
            I => buf_dds0_3
        );

    \I__8015\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40041\
        );

    \I__8014\ : CascadeMux
    port map (
            O => \N__40044\,
            I => \N__40038\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__40041\,
            I => \N__40035\
        );

    \I__8012\ : InMux
    port map (
            O => \N__40038\,
            I => \N__40032\
        );

    \I__8011\ : Span4Mux_v
    port map (
            O => \N__40035\,
            I => \N__40027\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__40032\,
            I => \N__40027\
        );

    \I__8009\ : Odrv4
    port map (
            O => \N__40027\,
            I => tmp_buf_15
        );

    \I__8008\ : IoInMux
    port map (
            O => \N__40024\,
            I => \N__40021\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__40021\,
            I => \N__40018\
        );

    \I__8006\ : Span4Mux_s2_v
    port map (
            O => \N__40018\,
            I => \N__40015\
        );

    \I__8005\ : Span4Mux_v
    port map (
            O => \N__40015\,
            I => \N__40012\
        );

    \I__8004\ : Sp12to4
    port map (
            O => \N__40012\,
            I => \N__40008\
        );

    \I__8003\ : InMux
    port map (
            O => \N__40011\,
            I => \N__40005\
        );

    \I__8002\ : Odrv12
    port map (
            O => \N__40008\,
            I => \DDS_MOSI\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__40005\,
            I => \DDS_MOSI\
        );

    \I__8000\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39997\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__39997\,
            I => \comm_spi.n24016\
        );

    \I__7998\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39991\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__39991\,
            I => \comm_spi.n15326\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__39988\,
            I => \comm_spi.n24016_cascade_\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__39985\,
            I => \n14_adj_1610_cascade_\
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__39982\,
            I => \N__39978\
        );

    \I__7993\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39975\
        );

    \I__7992\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39972\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__39975\,
            I => \N__39969\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__39972\,
            I => acadc_skipcnt_0
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__39969\,
            I => acadc_skipcnt_0
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__39964\,
            I => \N__39961\
        );

    \I__7987\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39958\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__39958\,
            I => \N__39954\
        );

    \I__7985\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39951\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__39954\,
            I => \N__39948\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__39951\,
            I => acadc_skipcnt_6
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__39948\,
            I => acadc_skipcnt_6
        );

    \I__7981\ : IoInMux
    port map (
            O => \N__39943\,
            I => \N__39940\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__39940\,
            I => \N__39937\
        );

    \I__7979\ : Span4Mux_s0_v
    port map (
            O => \N__39937\,
            I => \N__39934\
        );

    \I__7978\ : Span4Mux_v
    port map (
            O => \N__39934\,
            I => \N__39931\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__39931\,
            I => \N__39928\
        );

    \I__7976\ : Sp12to4
    port map (
            O => \N__39928\,
            I => \N__39923\
        );

    \I__7975\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39920\
        );

    \I__7974\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39917\
        );

    \I__7973\ : Odrv12
    port map (
            O => \N__39923\,
            I => \SELIRNG0\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__39920\,
            I => \SELIRNG0\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__39917\,
            I => \SELIRNG0\
        );

    \I__7970\ : InMux
    port map (
            O => \N__39910\,
            I => \N__39905\
        );

    \I__7969\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39902\
        );

    \I__7968\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39899\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__39905\,
            I => \acadc_skipCount_10\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__39902\,
            I => \acadc_skipCount_10\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__39899\,
            I => \acadc_skipCount_10\
        );

    \I__7964\ : IoInMux
    port map (
            O => \N__39892\,
            I => \N__39889\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__39889\,
            I => \N__39886\
        );

    \I__7962\ : Span4Mux_s0_h
    port map (
            O => \N__39886\,
            I => \N__39883\
        );

    \I__7961\ : Sp12to4
    port map (
            O => \N__39883\,
            I => \N__39880\
        );

    \I__7960\ : Span12Mux_v
    port map (
            O => \N__39880\,
            I => \N__39876\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__39879\,
            I => \N__39872\
        );

    \I__7958\ : Span12Mux_h
    port map (
            O => \N__39876\,
            I => \N__39869\
        );

    \I__7957\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39866\
        );

    \I__7956\ : InMux
    port map (
            O => \N__39872\,
            I => \N__39863\
        );

    \I__7955\ : Odrv12
    port map (
            O => \N__39869\,
            I => \VDC_RNG0\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__39866\,
            I => \VDC_RNG0\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__39863\,
            I => \VDC_RNG0\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__39856\,
            I => \N__39851\
        );

    \I__7951\ : CascadeMux
    port map (
            O => \N__39855\,
            I => \N__39848\
        );

    \I__7950\ : InMux
    port map (
            O => \N__39854\,
            I => \N__39845\
        );

    \I__7949\ : InMux
    port map (
            O => \N__39851\,
            I => \N__39840\
        );

    \I__7948\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39840\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__39845\,
            I => \acadc_skipCount_12\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__39840\,
            I => \acadc_skipCount_12\
        );

    \I__7945\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39832\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__39832\,
            I => \N__39829\
        );

    \I__7943\ : Span4Mux_v
    port map (
            O => \N__39829\,
            I => \N__39826\
        );

    \I__7942\ : Span4Mux_h
    port map (
            O => \N__39826\,
            I => \N__39823\
        );

    \I__7941\ : Odrv4
    port map (
            O => \N__39823\,
            I => n23_adj_1783
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__39820\,
            I => \N__39813\
        );

    \I__7939\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39801\
        );

    \I__7938\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39801\
        );

    \I__7937\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39794\
        );

    \I__7936\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39785\
        );

    \I__7935\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39785\
        );

    \I__7934\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39785\
        );

    \I__7933\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39785\
        );

    \I__7932\ : InMux
    port map (
            O => \N__39810\,
            I => \N__39782\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__39809\,
            I => \N__39777\
        );

    \I__7930\ : CascadeMux
    port map (
            O => \N__39808\,
            I => \N__39769\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__39807\,
            I => \N__39759\
        );

    \I__7928\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39755\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__39801\,
            I => \N__39750\
        );

    \I__7926\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39747\
        );

    \I__7925\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39738\
        );

    \I__7924\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39738\
        );

    \I__7923\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39738\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39733\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__39785\,
            I => \N__39733\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39729\
        );

    \I__7919\ : InMux
    port map (
            O => \N__39781\,
            I => \N__39725\
        );

    \I__7918\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39716\
        );

    \I__7917\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39716\
        );

    \I__7916\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39716\
        );

    \I__7915\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39716\
        );

    \I__7914\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39704\
        );

    \I__7913\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39704\
        );

    \I__7912\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39704\
        );

    \I__7911\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39701\
        );

    \I__7910\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39690\
        );

    \I__7909\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39690\
        );

    \I__7908\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39690\
        );

    \I__7907\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39690\
        );

    \I__7906\ : InMux
    port map (
            O => \N__39764\,
            I => \N__39690\
        );

    \I__7905\ : InMux
    port map (
            O => \N__39763\,
            I => \N__39685\
        );

    \I__7904\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39685\
        );

    \I__7903\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39682\
        );

    \I__7902\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39679\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39676\
        );

    \I__7900\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39672\
        );

    \I__7899\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39669\
        );

    \I__7898\ : Span4Mux_v
    port map (
            O => \N__39750\,
            I => \N__39664\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39664\
        );

    \I__7896\ : InMux
    port map (
            O => \N__39746\,
            I => \N__39659\
        );

    \I__7895\ : InMux
    port map (
            O => \N__39745\,
            I => \N__39659\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__39738\,
            I => \N__39656\
        );

    \I__7893\ : Span4Mux_v
    port map (
            O => \N__39733\,
            I => \N__39653\
        );

    \I__7892\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39648\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__39729\,
            I => \N__39645\
        );

    \I__7890\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39642\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__39725\,
            I => \N__39637\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__39716\,
            I => \N__39637\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__39715\,
            I => \N__39633\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__39714\,
            I => \N__39627\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__39713\,
            I => \N__39624\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__39712\,
            I => \N__39614\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__39711\,
            I => \N__39611\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39605\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__39701\,
            I => \N__39598\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__39690\,
            I => \N__39598\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__39685\,
            I => \N__39598\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__39682\,
            I => \N__39593\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39593\
        );

    \I__7876\ : Span4Mux_v
    port map (
            O => \N__39676\,
            I => \N__39590\
        );

    \I__7875\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39587\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39580\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__39669\,
            I => \N__39580\
        );

    \I__7872\ : Span4Mux_h
    port map (
            O => \N__39664\,
            I => \N__39580\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__39659\,
            I => \N__39573\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__39656\,
            I => \N__39573\
        );

    \I__7869\ : Span4Mux_v
    port map (
            O => \N__39653\,
            I => \N__39573\
        );

    \I__7868\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39568\
        );

    \I__7867\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39568\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__39648\,
            I => \N__39565\
        );

    \I__7865\ : Span4Mux_h
    port map (
            O => \N__39645\,
            I => \N__39562\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39557\
        );

    \I__7863\ : Span4Mux_v
    port map (
            O => \N__39637\,
            I => \N__39557\
        );

    \I__7862\ : InMux
    port map (
            O => \N__39636\,
            I => \N__39545\
        );

    \I__7861\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39542\
        );

    \I__7860\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39537\
        );

    \I__7859\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39537\
        );

    \I__7858\ : InMux
    port map (
            O => \N__39630\,
            I => \N__39534\
        );

    \I__7857\ : InMux
    port map (
            O => \N__39627\,
            I => \N__39523\
        );

    \I__7856\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39523\
        );

    \I__7855\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39523\
        );

    \I__7854\ : InMux
    port map (
            O => \N__39622\,
            I => \N__39523\
        );

    \I__7853\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39523\
        );

    \I__7852\ : InMux
    port map (
            O => \N__39620\,
            I => \N__39520\
        );

    \I__7851\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39513\
        );

    \I__7850\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39513\
        );

    \I__7849\ : InMux
    port map (
            O => \N__39617\,
            I => \N__39513\
        );

    \I__7848\ : InMux
    port map (
            O => \N__39614\,
            I => \N__39502\
        );

    \I__7847\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39502\
        );

    \I__7846\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39502\
        );

    \I__7845\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39502\
        );

    \I__7844\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39502\
        );

    \I__7843\ : Span4Mux_h
    port map (
            O => \N__39605\,
            I => \N__39499\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__39598\,
            I => \N__39496\
        );

    \I__7841\ : Span12Mux_h
    port map (
            O => \N__39593\,
            I => \N__39493\
        );

    \I__7840\ : Span4Mux_h
    port map (
            O => \N__39590\,
            I => \N__39490\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__39587\,
            I => \N__39483\
        );

    \I__7838\ : Span4Mux_v
    port map (
            O => \N__39580\,
            I => \N__39483\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__39573\,
            I => \N__39483\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__39568\,
            I => \N__39474\
        );

    \I__7835\ : Span4Mux_h
    port map (
            O => \N__39565\,
            I => \N__39474\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__39562\,
            I => \N__39474\
        );

    \I__7833\ : Span4Mux_h
    port map (
            O => \N__39557\,
            I => \N__39474\
        );

    \I__7832\ : InMux
    port map (
            O => \N__39556\,
            I => \N__39465\
        );

    \I__7831\ : InMux
    port map (
            O => \N__39555\,
            I => \N__39465\
        );

    \I__7830\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39465\
        );

    \I__7829\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39465\
        );

    \I__7828\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39454\
        );

    \I__7827\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39454\
        );

    \I__7826\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39454\
        );

    \I__7825\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39454\
        );

    \I__7824\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39454\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__39545\,
            I => adc_state_0
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__39542\,
            I => adc_state_0
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__39537\,
            I => adc_state_0
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__39534\,
            I => adc_state_0
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__39523\,
            I => adc_state_0
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__39520\,
            I => adc_state_0
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__39513\,
            I => adc_state_0
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__39502\,
            I => adc_state_0
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__39499\,
            I => adc_state_0
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__39496\,
            I => adc_state_0
        );

    \I__7813\ : Odrv12
    port map (
            O => \N__39493\,
            I => adc_state_0
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__39490\,
            I => adc_state_0
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__39483\,
            I => adc_state_0
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__39474\,
            I => adc_state_0
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__39465\,
            I => adc_state_0
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__39454\,
            I => adc_state_0
        );

    \I__7807\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39415\
        );

    \I__7806\ : InMux
    port map (
            O => \N__39420\,
            I => \N__39410\
        );

    \I__7805\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39410\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__39418\,
            I => \N__39407\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__39415\,
            I => \N__39395\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__39410\,
            I => \N__39392\
        );

    \I__7801\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39387\
        );

    \I__7800\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39387\
        );

    \I__7799\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39382\
        );

    \I__7798\ : InMux
    port map (
            O => \N__39404\,
            I => \N__39379\
        );

    \I__7797\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39372\
        );

    \I__7796\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39372\
        );

    \I__7795\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39365\
        );

    \I__7794\ : InMux
    port map (
            O => \N__39400\,
            I => \N__39365\
        );

    \I__7793\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39362\
        );

    \I__7792\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39357\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__39395\,
            I => \N__39352\
        );

    \I__7790\ : Span4Mux_h
    port map (
            O => \N__39392\,
            I => \N__39352\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__39387\,
            I => \N__39348\
        );

    \I__7788\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39345\
        );

    \I__7787\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39342\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__39382\,
            I => \N__39338\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__39379\,
            I => \N__39335\
        );

    \I__7784\ : InMux
    port map (
            O => \N__39378\,
            I => \N__39329\
        );

    \I__7783\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39329\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39326\
        );

    \I__7781\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39321\
        );

    \I__7780\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39321\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39318\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__39362\,
            I => \N__39315\
        );

    \I__7777\ : InMux
    port map (
            O => \N__39361\,
            I => \N__39310\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39310\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39305\
        );

    \I__7774\ : Span4Mux_v
    port map (
            O => \N__39352\,
            I => \N__39305\
        );

    \I__7773\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39302\
        );

    \I__7772\ : Span4Mux_h
    port map (
            O => \N__39348\,
            I => \N__39297\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39297\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__39342\,
            I => \N__39294\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39291\
        );

    \I__7768\ : Span4Mux_h
    port map (
            O => \N__39338\,
            I => \N__39286\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__39335\,
            I => \N__39286\
        );

    \I__7766\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39283\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__39329\,
            I => \N__39274\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__39326\,
            I => \N__39274\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__39321\,
            I => \N__39274\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__39318\,
            I => \N__39274\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__39315\,
            I => \N__39271\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39266\
        );

    \I__7759\ : Span4Mux_v
    port map (
            O => \N__39305\,
            I => \N__39266\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__39302\,
            I => \N__39263\
        );

    \I__7757\ : Span4Mux_v
    port map (
            O => \N__39297\,
            I => \N__39260\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__39294\,
            I => \N__39257\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__39291\,
            I => \N__39252\
        );

    \I__7754\ : Span4Mux_v
    port map (
            O => \N__39286\,
            I => \N__39252\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39283\,
            I => \N__39249\
        );

    \I__7752\ : Span4Mux_h
    port map (
            O => \N__39274\,
            I => \N__39246\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__39271\,
            I => \N__39241\
        );

    \I__7750\ : Span4Mux_h
    port map (
            O => \N__39266\,
            I => \N__39241\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__39263\,
            I => \N__39232\
        );

    \I__7748\ : Span4Mux_h
    port map (
            O => \N__39260\,
            I => \N__39232\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__39257\,
            I => \N__39232\
        );

    \I__7746\ : Span4Mux_h
    port map (
            O => \N__39252\,
            I => \N__39232\
        );

    \I__7745\ : Odrv4
    port map (
            O => \N__39249\,
            I => n21951
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__39246\,
            I => n21951
        );

    \I__7743\ : Odrv4
    port map (
            O => \N__39241\,
            I => n21951
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__39232\,
            I => n21951
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__7740\ : InMux
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__39217\,
            I => \N__39213\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__39216\,
            I => \N__39210\
        );

    \I__7737\ : Span12Mux_h
    port map (
            O => \N__39213\,
            I => \N__39206\
        );

    \I__7736\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39201\
        );

    \I__7735\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39201\
        );

    \I__7734\ : Odrv12
    port map (
            O => \N__39206\,
            I => cmd_rdadctmp_17
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39201\,
            I => cmd_rdadctmp_17
        );

    \I__7732\ : InMux
    port map (
            O => \N__39196\,
            I => \N__39193\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__39193\,
            I => \N__39188\
        );

    \I__7730\ : InMux
    port map (
            O => \N__39192\,
            I => \N__39183\
        );

    \I__7729\ : InMux
    port map (
            O => \N__39191\,
            I => \N__39183\
        );

    \I__7728\ : Odrv4
    port map (
            O => \N__39188\,
            I => req_data_cnt_10
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__39183\,
            I => req_data_cnt_10
        );

    \I__7726\ : SRMux
    port map (
            O => \N__39178\,
            I => \N__39174\
        );

    \I__7725\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39167\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__39174\,
            I => \N__39164\
        );

    \I__7723\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39161\
        );

    \I__7722\ : SRMux
    port map (
            O => \N__39172\,
            I => \N__39158\
        );

    \I__7721\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39155\
        );

    \I__7720\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39152\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__39167\,
            I => \N__39149\
        );

    \I__7718\ : Span4Mux_v
    port map (
            O => \N__39164\,
            I => \N__39145\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__39161\,
            I => \N__39142\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__39158\,
            I => \N__39137\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__39155\,
            I => \N__39137\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__39152\,
            I => \N__39134\
        );

    \I__7713\ : Span12Mux_s10_v
    port map (
            O => \N__39149\,
            I => \N__39127\
        );

    \I__7712\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39124\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__39145\,
            I => \N__39119\
        );

    \I__7710\ : Span4Mux_v
    port map (
            O => \N__39142\,
            I => \N__39119\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__39137\,
            I => \N__39116\
        );

    \I__7708\ : Span12Mux_h
    port map (
            O => \N__39134\,
            I => \N__39113\
        );

    \I__7707\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39110\
        );

    \I__7706\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39105\
        );

    \I__7705\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39105\
        );

    \I__7704\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39102\
        );

    \I__7703\ : Odrv12
    port map (
            O => \N__39127\,
            I => acadc_rst
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__39124\,
            I => acadc_rst
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__39119\,
            I => acadc_rst
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__39116\,
            I => acadc_rst
        );

    \I__7699\ : Odrv12
    port map (
            O => \N__39113\,
            I => acadc_rst
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__39110\,
            I => acadc_rst
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__39105\,
            I => acadc_rst
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__39102\,
            I => acadc_rst
        );

    \I__7695\ : CascadeMux
    port map (
            O => \N__39085\,
            I => \N__39082\
        );

    \I__7694\ : CascadeBuf
    port map (
            O => \N__39082\,
            I => \N__39079\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__39079\,
            I => \N__39076\
        );

    \I__7692\ : CascadeBuf
    port map (
            O => \N__39076\,
            I => \N__39073\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__39073\,
            I => \N__39070\
        );

    \I__7690\ : CascadeBuf
    port map (
            O => \N__39070\,
            I => \N__39067\
        );

    \I__7689\ : CascadeMux
    port map (
            O => \N__39067\,
            I => \N__39064\
        );

    \I__7688\ : CascadeBuf
    port map (
            O => \N__39064\,
            I => \N__39061\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__39061\,
            I => \N__39058\
        );

    \I__7686\ : CascadeBuf
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__7685\ : CascadeMux
    port map (
            O => \N__39055\,
            I => \N__39052\
        );

    \I__7684\ : CascadeBuf
    port map (
            O => \N__39052\,
            I => \N__39049\
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__39049\,
            I => \N__39046\
        );

    \I__7682\ : CascadeBuf
    port map (
            O => \N__39046\,
            I => \N__39042\
        );

    \I__7681\ : CascadeMux
    port map (
            O => \N__39045\,
            I => \N__39039\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__39042\,
            I => \N__39036\
        );

    \I__7679\ : CascadeBuf
    port map (
            O => \N__39039\,
            I => \N__39033\
        );

    \I__7678\ : CascadeBuf
    port map (
            O => \N__39036\,
            I => \N__39030\
        );

    \I__7677\ : CascadeMux
    port map (
            O => \N__39033\,
            I => \N__39027\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__39030\,
            I => \N__39024\
        );

    \I__7675\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39021\
        );

    \I__7674\ : CascadeBuf
    port map (
            O => \N__39024\,
            I => \N__39018\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__39021\,
            I => \N__39015\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__39018\,
            I => \N__39012\
        );

    \I__7671\ : Span4Mux_v
    port map (
            O => \N__39015\,
            I => \N__39009\
        );

    \I__7670\ : InMux
    port map (
            O => \N__39012\,
            I => \N__39006\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__39009\,
            I => \N__39003\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__39006\,
            I => \N__39000\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__39003\,
            I => \N__38997\
        );

    \I__7666\ : Span4Mux_v
    port map (
            O => \N__39000\,
            I => \N__38994\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__38997\,
            I => \N__38991\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__38994\,
            I => \N__38988\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__38991\,
            I => \data_index_9_N_236_3\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__38988\,
            I => \data_index_9_N_236_3\
        );

    \I__7661\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38980\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__38980\,
            I => \N__38976\
        );

    \I__7659\ : InMux
    port map (
            O => \N__38979\,
            I => \N__38973\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__38976\,
            I => \N__38970\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__38973\,
            I => acadc_skipcnt_7
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__38970\,
            I => acadc_skipcnt_7
        );

    \I__7655\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38958\
        );

    \I__7653\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38955\
        );

    \I__7652\ : Span4Mux_h
    port map (
            O => \N__38958\,
            I => \N__38952\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__38955\,
            I => acadc_skipcnt_2
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__38952\,
            I => acadc_skipcnt_2
        );

    \I__7649\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38944\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__38944\,
            I => \N__38940\
        );

    \I__7647\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38937\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__38940\,
            I => \N__38934\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__38937\,
            I => acadc_skipcnt_12
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__38934\,
            I => acadc_skipcnt_12
        );

    \I__7643\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38926\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38922\
        );

    \I__7641\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38919\
        );

    \I__7640\ : Span4Mux_h
    port map (
            O => \N__38922\,
            I => \N__38916\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__38919\,
            I => acadc_skipcnt_10
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__38916\,
            I => acadc_skipcnt_10
        );

    \I__7637\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38905\
        );

    \I__7635\ : Odrv4
    port map (
            O => \N__38905\,
            I => n23_adj_1514
        );

    \I__7634\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38899\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__38899\,
            I => n24_adj_1513
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__38896\,
            I => \n21_cascade_\
        );

    \I__7631\ : InMux
    port map (
            O => \N__38893\,
            I => \N__38890\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__38890\,
            I => n22
        );

    \I__7629\ : InMux
    port map (
            O => \N__38887\,
            I => n20656
        );

    \I__7628\ : InMux
    port map (
            O => \N__38884\,
            I => n20657
        );

    \I__7627\ : InMux
    port map (
            O => \N__38881\,
            I => n20658
        );

    \I__7626\ : InMux
    port map (
            O => \N__38878\,
            I => \bfn_13_16_0_\
        );

    \I__7625\ : InMux
    port map (
            O => \N__38875\,
            I => n20660
        );

    \I__7624\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38868\
        );

    \I__7623\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38863\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__38868\,
            I => \N__38860\
        );

    \I__7621\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38857\
        );

    \I__7620\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38854\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__38863\,
            I => \N__38851\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__38860\,
            I => \N__38846\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__38857\,
            I => \N__38846\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__38854\,
            I => eis_stop
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__38851\,
            I => eis_stop
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__38846\,
            I => eis_stop
        );

    \I__7613\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38836\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__38836\,
            I => \N__38832\
        );

    \I__7611\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38829\
        );

    \I__7610\ : Span4Mux_h
    port map (
            O => \N__38832\,
            I => \N__38826\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__38829\,
            I => acadc_skipcnt_13
        );

    \I__7608\ : Odrv4
    port map (
            O => \N__38826\,
            I => acadc_skipcnt_13
        );

    \I__7607\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38818\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__38818\,
            I => \N__38813\
        );

    \I__7605\ : InMux
    port map (
            O => \N__38817\,
            I => \N__38808\
        );

    \I__7604\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38808\
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__38813\,
            I => \acadc_skipCount_13\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__38808\,
            I => \acadc_skipCount_13\
        );

    \I__7601\ : IoInMux
    port map (
            O => \N__38803\,
            I => \N__38800\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__7599\ : Span12Mux_s3_h
    port map (
            O => \N__38797\,
            I => \N__38794\
        );

    \I__7598\ : Span12Mux_h
    port map (
            O => \N__38794\,
            I => \N__38789\
        );

    \I__7597\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38786\
        );

    \I__7596\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38783\
        );

    \I__7595\ : Odrv12
    port map (
            O => \N__38789\,
            I => \VAC_OSR0\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__38786\,
            I => \VAC_OSR0\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__38783\,
            I => \VAC_OSR0\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__38776\,
            I => \N__38769\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__38775\,
            I => \N__38766\
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__38774\,
            I => \N__38763\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__38773\,
            I => \N__38760\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__38772\,
            I => \N__38754\
        );

    \I__7587\ : InMux
    port map (
            O => \N__38769\,
            I => \N__38747\
        );

    \I__7586\ : InMux
    port map (
            O => \N__38766\,
            I => \N__38747\
        );

    \I__7585\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38747\
        );

    \I__7584\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38744\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__38759\,
            I => \N__38741\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__38758\,
            I => \N__38738\
        );

    \I__7581\ : InMux
    port map (
            O => \N__38757\,
            I => \N__38733\
        );

    \I__7580\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38733\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__38747\,
            I => \N__38730\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__38744\,
            I => \N__38727\
        );

    \I__7577\ : InMux
    port map (
            O => \N__38741\,
            I => \N__38722\
        );

    \I__7576\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38722\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__38733\,
            I => \N__38719\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__38730\,
            I => \N__38712\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__38727\,
            I => \N__38712\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__38722\,
            I => \N__38712\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__38719\,
            I => n40
        );

    \I__7570\ : Odrv4
    port map (
            O => \N__38712\,
            I => n40
        );

    \I__7569\ : InMux
    port map (
            O => \N__38707\,
            I => \N__38704\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__38704\,
            I => \N__38701\
        );

    \I__7567\ : Odrv4
    port map (
            O => \N__38701\,
            I => n24_adj_1505
        );

    \I__7566\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38695\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__38695\,
            I => \N__38691\
        );

    \I__7564\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38687\
        );

    \I__7563\ : Span4Mux_h
    port map (
            O => \N__38691\,
            I => \N__38684\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__38690\,
            I => \N__38681\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38676\
        );

    \I__7560\ : Span4Mux_h
    port map (
            O => \N__38684\,
            I => \N__38676\
        );

    \I__7559\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38673\
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__38676\,
            I => req_data_cnt_12
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__38673\,
            I => req_data_cnt_12
        );

    \I__7556\ : IoInMux
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__38665\,
            I => \N__38662\
        );

    \I__7554\ : Span4Mux_s2_h
    port map (
            O => \N__38662\,
            I => \N__38658\
        );

    \I__7553\ : InMux
    port map (
            O => \N__38661\,
            I => \N__38654\
        );

    \I__7552\ : Sp12to4
    port map (
            O => \N__38658\,
            I => \N__38651\
        );

    \I__7551\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38648\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38645\
        );

    \I__7549\ : Span12Mux_v
    port map (
            O => \N__38651\,
            I => \N__38642\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__38648\,
            I => \N__38639\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__38645\,
            I => \N__38636\
        );

    \I__7546\ : Span12Mux_h
    port map (
            O => \N__38642\,
            I => \N__38633\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__38639\,
            I => \N__38628\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__38636\,
            I => \N__38628\
        );

    \I__7543\ : Odrv12
    port map (
            O => \N__38633\,
            I => \VAC_OSR1\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__38628\,
            I => \VAC_OSR1\
        );

    \I__7541\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38620\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__38620\,
            I => \N__38616\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__38619\,
            I => \N__38613\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__38616\,
            I => \N__38610\
        );

    \I__7537\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38607\
        );

    \I__7536\ : Sp12to4
    port map (
            O => \N__38610\,
            I => \N__38603\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__38607\,
            I => \N__38600\
        );

    \I__7534\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38597\
        );

    \I__7533\ : Span12Mux_h
    port map (
            O => \N__38603\,
            I => \N__38594\
        );

    \I__7532\ : Span4Mux_h
    port map (
            O => \N__38600\,
            I => \N__38591\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__38597\,
            I => buf_adcdata_iac_21
        );

    \I__7530\ : Odrv12
    port map (
            O => \N__38594\,
            I => buf_adcdata_iac_21
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__38591\,
            I => buf_adcdata_iac_21
        );

    \I__7528\ : InMux
    port map (
            O => \N__38584\,
            I => \N__38579\
        );

    \I__7527\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38576\
        );

    \I__7526\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38573\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38570\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__38576\,
            I => \N__38565\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__38573\,
            I => \N__38565\
        );

    \I__7522\ : Odrv12
    port map (
            O => \N__38570\,
            I => n9_adj_1600
        );

    \I__7521\ : Odrv4
    port map (
            O => \N__38565\,
            I => n9_adj_1600
        );

    \I__7520\ : InMux
    port map (
            O => \N__38560\,
            I => \bfn_13_15_0_\
        );

    \I__7519\ : InMux
    port map (
            O => \N__38557\,
            I => n20652
        );

    \I__7518\ : InMux
    port map (
            O => \N__38554\,
            I => n20653
        );

    \I__7517\ : InMux
    port map (
            O => \N__38551\,
            I => n20654
        );

    \I__7516\ : InMux
    port map (
            O => \N__38548\,
            I => n20655
        );

    \I__7515\ : CascadeMux
    port map (
            O => \N__38545\,
            I => \n23450_cascade_\
        );

    \I__7514\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38539\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__38539\,
            I => \N__38536\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__38536\,
            I => \N__38533\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__38533\,
            I => n23327
        );

    \I__7510\ : InMux
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__38527\,
            I => \N__38524\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__38524\,
            I => n23453
        );

    \I__7507\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__38515\,
            I => n112_adj_1583
        );

    \I__7504\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__38509\,
            I => \N__38506\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__38506\,
            I => \N__38503\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__38503\,
            I => n23522
        );

    \I__7500\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38497\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__38497\,
            I => n22267
        );

    \I__7498\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38491\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__38491\,
            I => n112_adj_1797
        );

    \I__7496\ : CascadeMux
    port map (
            O => \N__38488\,
            I => \N__38485\
        );

    \I__7495\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38482\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__38479\,
            I => \comm_buf_0_7_N_543_2\
        );

    \I__7492\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38469\
        );

    \I__7490\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38466\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__38469\,
            I => \N__38463\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__38466\,
            I => comm_test_buf_24_16
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__38463\,
            I => comm_test_buf_24_16
        );

    \I__7486\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38455\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__38455\,
            I => n111_adj_1584
        );

    \I__7484\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38449\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__38449\,
            I => \N__38446\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__38446\,
            I => n20_adj_1804
        );

    \I__7481\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38440\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__38440\,
            I => \N__38437\
        );

    \I__7479\ : Span4Mux_v
    port map (
            O => \N__38437\,
            I => \N__38433\
        );

    \I__7478\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38430\
        );

    \I__7477\ : Odrv4
    port map (
            O => \N__38433\,
            I => \comm_spi.n15338\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__38430\,
            I => \comm_spi.n15338\
        );

    \I__7475\ : SRMux
    port map (
            O => \N__38425\,
            I => \N__38422\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__38422\,
            I => \N__38419\
        );

    \I__7473\ : Odrv4
    port map (
            O => \N__38419\,
            I => n15496
        );

    \I__7472\ : CascadeMux
    port map (
            O => \N__38416\,
            I => \N__38413\
        );

    \I__7471\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38410\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__38410\,
            I => \N__38407\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__38407\,
            I => \N__38404\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__38404\,
            I => \N__38401\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__38401\,
            I => buf_data_iac_16
        );

    \I__7466\ : CascadeMux
    port map (
            O => \N__38398\,
            I => \n22270_cascade_\
        );

    \I__7465\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38388\
        );

    \I__7463\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38385\
        );

    \I__7462\ : Span4Mux_h
    port map (
            O => \N__38388\,
            I => \N__38382\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__38385\,
            I => comm_test_buf_24_9
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__38382\,
            I => comm_test_buf_24_9
        );

    \I__7459\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38374\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__38374\,
            I => \comm_buf_0_7_N_543_0\
        );

    \I__7457\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38368\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__38368\,
            I => \N__38364\
        );

    \I__7455\ : InMux
    port map (
            O => \N__38367\,
            I => \N__38361\
        );

    \I__7454\ : Span4Mux_v
    port map (
            O => \N__38364\,
            I => \N__38358\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__38361\,
            I => comm_test_buf_24_18
        );

    \I__7452\ : Odrv4
    port map (
            O => \N__38358\,
            I => comm_test_buf_24_18
        );

    \I__7451\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38348\
        );

    \I__7450\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38345\
        );

    \I__7449\ : InMux
    port map (
            O => \N__38351\,
            I => \N__38342\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__38348\,
            I => \N__38339\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__38345\,
            I => \N__38334\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__38342\,
            I => \N__38334\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__38339\,
            I => comm_test_buf_24_7
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__38334\,
            I => comm_test_buf_24_7
        );

    \I__7443\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38326\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__7441\ : Span4Mux_h
    port map (
            O => \N__38323\,
            I => \N__38319\
        );

    \I__7440\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38316\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__38319\,
            I => comm_test_buf_24_15
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__38316\,
            I => comm_test_buf_24_15
        );

    \I__7437\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__38308\,
            I => \N__38304\
        );

    \I__7435\ : InMux
    port map (
            O => \N__38307\,
            I => \N__38301\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__38304\,
            I => \N__38298\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__38301\,
            I => \N__38294\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__38298\,
            I => \N__38291\
        );

    \I__7431\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38288\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__38294\,
            I => \N__38285\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__38291\,
            I => comm_buf_2_1
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__38288\,
            I => comm_buf_2_1
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__38285\,
            I => comm_buf_2_1
        );

    \I__7426\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__38272\,
            I => \N__38269\
        );

    \I__7423\ : Odrv4
    port map (
            O => \N__38269\,
            I => n13201
        );

    \I__7422\ : InMux
    port map (
            O => \N__38266\,
            I => \N__38263\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__38263\,
            I => \N__38260\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__38260\,
            I => \N__38257\
        );

    \I__7419\ : Sp12to4
    port map (
            O => \N__38257\,
            I => \N__38253\
        );

    \I__7418\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38250\
        );

    \I__7417\ : Odrv12
    port map (
            O => \N__38253\,
            I => \buf_readRTD_9\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__38250\,
            I => \buf_readRTD_9\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__38245\,
            I => \N__38242\
        );

    \I__7414\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38239\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38234\
        );

    \I__7412\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38230\
        );

    \I__7411\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38227\
        );

    \I__7410\ : Span4Mux_v
    port map (
            O => \N__38234\,
            I => \N__38224\
        );

    \I__7409\ : InMux
    port map (
            O => \N__38233\,
            I => \N__38221\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__38230\,
            I => \N__38216\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38216\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__38224\,
            I => \N__38212\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__38221\,
            I => \N__38209\
        );

    \I__7404\ : Span12Mux_v
    port map (
            O => \N__38216\,
            I => \N__38206\
        );

    \I__7403\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38203\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__38212\,
            I => \N__38198\
        );

    \I__7401\ : Span4Mux_v
    port map (
            O => \N__38209\,
            I => \N__38198\
        );

    \I__7400\ : Odrv12
    port map (
            O => \N__38206\,
            I => \buf_cfgRTD_1\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__38203\,
            I => \buf_cfgRTD_1\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__38198\,
            I => \buf_cfgRTD_1\
        );

    \I__7397\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38188\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__7395\ : Span4Mux_v
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__38182\,
            I => \N__38178\
        );

    \I__7393\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38175\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__38178\,
            I => \comm_spi.n15337\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__38175\,
            I => \comm_spi.n15337\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__38170\,
            I => \N__38167\
        );

    \I__7389\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N__38161\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__38161\,
            I => \N__38157\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__38160\,
            I => \N__38154\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__38157\,
            I => \N__38151\
        );

    \I__7384\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38148\
        );

    \I__7383\ : Sp12to4
    port map (
            O => \N__38151\,
            I => \N__38145\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__38148\,
            I => cmd_rdadctmp_7
        );

    \I__7381\ : Odrv12
    port map (
            O => \N__38145\,
            I => cmd_rdadctmp_7
        );

    \I__7380\ : InMux
    port map (
            O => \N__38140\,
            I => \N__38136\
        );

    \I__7379\ : InMux
    port map (
            O => \N__38139\,
            I => \N__38133\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__38136\,
            I => comm_buf_6_4
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__38133\,
            I => comm_buf_6_4
        );

    \I__7376\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__7374\ : Span4Mux_v
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__7373\ : Span4Mux_h
    port map (
            O => \N__38119\,
            I => \N__38114\
        );

    \I__7372\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38111\
        );

    \I__7371\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38108\
        );

    \I__7370\ : Span4Mux_v
    port map (
            O => \N__38114\,
            I => \N__38105\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__38111\,
            I => cmd_rdadctmp_8
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__38108\,
            I => cmd_rdadctmp_8
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__38105\,
            I => cmd_rdadctmp_8
        );

    \I__7366\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38094\
        );

    \I__7365\ : CascadeMux
    port map (
            O => \N__38097\,
            I => \N__38091\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38094\,
            I => \N__38088\
        );

    \I__7363\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38084\
        );

    \I__7362\ : Span12Mux_v
    port map (
            O => \N__38088\,
            I => \N__38081\
        );

    \I__7361\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38078\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__38084\,
            I => buf_adcdata_iac_0
        );

    \I__7359\ : Odrv12
    port map (
            O => \N__38081\,
            I => buf_adcdata_iac_0
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__38078\,
            I => buf_adcdata_iac_0
        );

    \I__7357\ : InMux
    port map (
            O => \N__38071\,
            I => \N__38068\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__38068\,
            I => \N__38065\
        );

    \I__7355\ : Span4Mux_h
    port map (
            O => \N__38065\,
            I => \N__38062\
        );

    \I__7354\ : Span4Mux_v
    port map (
            O => \N__38062\,
            I => \N__38058\
        );

    \I__7353\ : InMux
    port map (
            O => \N__38061\,
            I => \N__38055\
        );

    \I__7352\ : Odrv4
    port map (
            O => \N__38058\,
            I => buf_adcdata_vdc_13
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__38055\,
            I => buf_adcdata_vdc_13
        );

    \I__7350\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38047\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__38044\,
            I => \N__38040\
        );

    \I__7347\ : InMux
    port map (
            O => \N__38043\,
            I => \N__38037\
        );

    \I__7346\ : Span4Mux_h
    port map (
            O => \N__38040\,
            I => \N__38033\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__38037\,
            I => \N__38030\
        );

    \I__7344\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38027\
        );

    \I__7343\ : Span4Mux_h
    port map (
            O => \N__38033\,
            I => \N__38022\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__38030\,
            I => \N__38022\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__38027\,
            I => buf_adcdata_vac_13
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__38022\,
            I => buf_adcdata_vac_13
        );

    \I__7339\ : InMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__38014\,
            I => \N__38011\
        );

    \I__7337\ : Span4Mux_v
    port map (
            O => \N__38011\,
            I => \N__38008\
        );

    \I__7336\ : Span4Mux_h
    port map (
            O => \N__38008\,
            I => \N__38005\
        );

    \I__7335\ : Span4Mux_h
    port map (
            O => \N__38005\,
            I => \N__38001\
        );

    \I__7334\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37998\
        );

    \I__7333\ : Odrv4
    port map (
            O => \N__38001\,
            I => \buf_readRTD_5\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__37998\,
            I => \buf_readRTD_5\
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__37993\,
            I => \n19_adj_1729_cascade_\
        );

    \I__7330\ : InMux
    port map (
            O => \N__37990\,
            I => \N__37986\
        );

    \I__7329\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37980\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__37983\,
            I => comm_buf_6_6
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__37980\,
            I => comm_buf_6_6
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__37975\,
            I => \n9_adj_1600_cascade_\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__37972\,
            I => \n6776_cascade_\
        );

    \I__7323\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37966\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__37963\,
            I => \N__37960\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__37960\,
            I => n18890
        );

    \I__7319\ : InMux
    port map (
            O => \N__37957\,
            I => \N__37954\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37951\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__37951\,
            I => \N__37948\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__37948\,
            I => n23390
        );

    \I__7315\ : CascadeMux
    port map (
            O => \N__37945\,
            I => \n1_adj_1674_cascade_\
        );

    \I__7314\ : InMux
    port map (
            O => \N__37942\,
            I => \N__37935\
        );

    \I__7313\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37935\
        );

    \I__7312\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37932\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__37935\,
            I => \N__37929\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37926\
        );

    \I__7309\ : Odrv12
    port map (
            O => \N__37929\,
            I => comm_tx_buf_1
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__37926\,
            I => comm_tx_buf_1
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__37921\,
            I => \N__37918\
        );

    \I__7306\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37915\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__37915\,
            I => \N__37912\
        );

    \I__7304\ : Odrv4
    port map (
            O => \N__37912\,
            I => n22341
        );

    \I__7303\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37906\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__37906\,
            I => n2_adj_1675
        );

    \I__7301\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37900\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__37900\,
            I => \N__37896\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__37899\,
            I => \N__37893\
        );

    \I__7298\ : Sp12to4
    port map (
            O => \N__37896\,
            I => \N__37890\
        );

    \I__7297\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37887\
        );

    \I__7296\ : Odrv12
    port map (
            O => \N__37890\,
            I => buf_adcdata_vdc_0
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__37887\,
            I => buf_adcdata_vdc_0
        );

    \I__7294\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37875\
        );

    \I__7292\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37871\
        );

    \I__7291\ : Span12Mux_s10_h
    port map (
            O => \N__37875\,
            I => \N__37868\
        );

    \I__7290\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37865\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__37871\,
            I => buf_adcdata_vac_0
        );

    \I__7288\ : Odrv12
    port map (
            O => \N__37868\,
            I => buf_adcdata_vac_0
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__37865\,
            I => buf_adcdata_vac_0
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__37858\,
            I => \n19_adj_1590_cascade_\
        );

    \I__7285\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37852\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__37852\,
            I => \N__37849\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__37846\,
            I => n22_adj_1589
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__37843\,
            I => \n21965_cascade_\
        );

    \I__7280\ : InMux
    port map (
            O => \N__37840\,
            I => \N__37833\
        );

    \I__7279\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37825\
        );

    \I__7278\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37825\
        );

    \I__7277\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37816\
        );

    \I__7276\ : InMux
    port map (
            O => \N__37836\,
            I => \N__37816\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__37833\,
            I => \N__37811\
        );

    \I__7274\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37807\
        );

    \I__7273\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37802\
        );

    \I__7272\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37802\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__37825\,
            I => \N__37797\
        );

    \I__7270\ : InMux
    port map (
            O => \N__37824\,
            I => \N__37786\
        );

    \I__7269\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37779\
        );

    \I__7268\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37779\
        );

    \I__7267\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37779\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37776\
        );

    \I__7265\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37773\
        );

    \I__7264\ : InMux
    port map (
            O => \N__37814\,
            I => \N__37769\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__37811\,
            I => \N__37766\
        );

    \I__7262\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37763\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37758\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__37802\,
            I => \N__37758\
        );

    \I__7259\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37755\
        );

    \I__7258\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37752\
        );

    \I__7257\ : Span4Mux_v
    port map (
            O => \N__37797\,
            I => \N__37749\
        );

    \I__7256\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37740\
        );

    \I__7255\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37737\
        );

    \I__7254\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37732\
        );

    \I__7253\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37732\
        );

    \I__7252\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37723\
        );

    \I__7251\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37723\
        );

    \I__7250\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37723\
        );

    \I__7249\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37723\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__37786\,
            I => \N__37718\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__37779\,
            I => \N__37718\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__37776\,
            I => \N__37713\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__37773\,
            I => \N__37713\
        );

    \I__7244\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37710\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__37769\,
            I => \N__37707\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__37766\,
            I => \N__37700\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37700\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__37758\,
            I => \N__37700\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__37755\,
            I => \N__37697\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__37752\,
            I => \N__37692\
        );

    \I__7237\ : Sp12to4
    port map (
            O => \N__37749\,
            I => \N__37692\
        );

    \I__7236\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37689\
        );

    \I__7235\ : InMux
    port map (
            O => \N__37747\,
            I => \N__37678\
        );

    \I__7234\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37678\
        );

    \I__7233\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37678\
        );

    \I__7232\ : InMux
    port map (
            O => \N__37744\,
            I => \N__37678\
        );

    \I__7231\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37678\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__37740\,
            I => \N__37671\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37671\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__37732\,
            I => \N__37671\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__37723\,
            I => \N__37668\
        );

    \I__7226\ : Span4Mux_v
    port map (
            O => \N__37718\,
            I => \N__37665\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__37713\,
            I => \N__37662\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__37710\,
            I => \N__37655\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__37707\,
            I => \N__37655\
        );

    \I__7222\ : Span4Mux_h
    port map (
            O => \N__37700\,
            I => \N__37655\
        );

    \I__7221\ : Sp12to4
    port map (
            O => \N__37697\,
            I => \N__37650\
        );

    \I__7220\ : Span12Mux_h
    port map (
            O => \N__37692\,
            I => \N__37650\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__37689\,
            I => n13746
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__37678\,
            I => n13746
        );

    \I__7217\ : Odrv12
    port map (
            O => \N__37671\,
            I => n13746
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__37668\,
            I => n13746
        );

    \I__7215\ : Odrv4
    port map (
            O => \N__37665\,
            I => n13746
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__37662\,
            I => n13746
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__37655\,
            I => n13746
        );

    \I__7212\ : Odrv12
    port map (
            O => \N__37650\,
            I => n13746
        );

    \I__7211\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37630\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__37630\,
            I => \N__37627\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__37627\,
            I => \N__37623\
        );

    \I__7208\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37620\
        );

    \I__7207\ : Sp12to4
    port map (
            O => \N__37623\,
            I => \N__37615\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37615\
        );

    \I__7205\ : Odrv12
    port map (
            O => \N__37615\,
            I => \comm_spi.n15323\
        );

    \I__7204\ : SRMux
    port map (
            O => \N__37612\,
            I => \N__37609\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__37609\,
            I => \N__37606\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__37606\,
            I => \comm_spi.data_tx_7__N_860\
        );

    \I__7201\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37600\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37595\
        );

    \I__7199\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37592\
        );

    \I__7198\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37589\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__37595\,
            I => \comm_spi.n24040\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__37592\,
            I => \comm_spi.n24040\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__37589\,
            I => \comm_spi.n24040\
        );

    \I__7194\ : SRMux
    port map (
            O => \N__37582\,
            I => \N__37579\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__37579\,
            I => \N__37576\
        );

    \I__7192\ : Odrv12
    port map (
            O => \N__37576\,
            I => \comm_spi.data_tx_7__N_880\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__37573\,
            I => \N__37570\
        );

    \I__7190\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37567\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37564\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__37564\,
            I => \N__37560\
        );

    \I__7187\ : InMux
    port map (
            O => \N__37563\,
            I => \N__37557\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__37560\,
            I => \N__37553\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37550\
        );

    \I__7184\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37547\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__37553\,
            I => \comm_spi.n24037\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__37550\,
            I => \comm_spi.n24037\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__37547\,
            I => \comm_spi.n24037\
        );

    \I__7180\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37537\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__37537\,
            I => \N__37534\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__37534\,
            I => \N__37530\
        );

    \I__7177\ : InMux
    port map (
            O => \N__37533\,
            I => \N__37527\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__37530\,
            I => \N__37522\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__37527\,
            I => \N__37522\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__37522\,
            I => \comm_spi.n15348\
        );

    \I__7173\ : InMux
    port map (
            O => \N__37519\,
            I => \N__37516\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37513\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__37513\,
            I => \N__37510\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__37510\,
            I => \N__37506\
        );

    \I__7169\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37503\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__37506\,
            I => \N__37500\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37497\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__37500\,
            I => \comm_spi.n15349\
        );

    \I__7165\ : Odrv12
    port map (
            O => \N__37497\,
            I => \comm_spi.n15349\
        );

    \I__7164\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37489\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__37489\,
            I => \comm_spi.n15335\
        );

    \I__7162\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37480\
        );

    \I__7161\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37480\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__37480\,
            I => buf_control_6
        );

    \I__7159\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37472\
        );

    \I__7158\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37467\
        );

    \I__7157\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37467\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__37472\,
            I => \acadc_skipCount_14\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__37467\,
            I => \acadc_skipCount_14\
        );

    \I__7154\ : CascadeMux
    port map (
            O => \N__37462\,
            I => \N__37459\
        );

    \I__7153\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37456\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__7151\ : Span12Mux_h
    port map (
            O => \N__37453\,
            I => \N__37450\
        );

    \I__7150\ : Odrv12
    port map (
            O => \N__37450\,
            I => n23_adj_1767
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__37447\,
            I => \N__37444\
        );

    \I__7148\ : InMux
    port map (
            O => \N__37444\,
            I => \N__37441\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__37441\,
            I => \SIG_DDS.tmp_buf_0\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__37438\,
            I => \N__37435\
        );

    \I__7145\ : InMux
    port map (
            O => \N__37435\,
            I => \N__37432\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__37432\,
            I => \N__37429\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__37429\,
            I => \N__37426\
        );

    \I__7142\ : Odrv4
    port map (
            O => \N__37426\,
            I => \SIG_DDS.tmp_buf_3\
        );

    \I__7141\ : CascadeMux
    port map (
            O => \N__37423\,
            I => \N__37420\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37420\,
            I => \N__37417\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__37417\,
            I => \SIG_DDS.tmp_buf_1\
        );

    \I__7138\ : CascadeMux
    port map (
            O => \N__37414\,
            I => \N__37411\
        );

    \I__7137\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37408\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__37408\,
            I => \SIG_DDS.tmp_buf_2\
        );

    \I__7135\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37398\
        );

    \I__7134\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__7133\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37395\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__37398\,
            I => \N__37389\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__37395\,
            I => \N__37386\
        );

    \I__7130\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37383\
        );

    \I__7129\ : InMux
    port map (
            O => \N__37393\,
            I => \N__37376\
        );

    \I__7128\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37376\
        );

    \I__7127\ : Span4Mux_h
    port map (
            O => \N__37389\,
            I => \N__37373\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__37386\,
            I => \N__37368\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__37383\,
            I => \N__37368\
        );

    \I__7124\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37365\
        );

    \I__7123\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37362\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37376\,
            I => n11979
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__37373\,
            I => n11979
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__37368\,
            I => n11979
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__37365\,
            I => n11979
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__37362\,
            I => n11979
        );

    \I__7117\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37348\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__37348\,
            I => \N__37344\
        );

    \I__7115\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37341\
        );

    \I__7114\ : Span4Mux_h
    port map (
            O => \N__37344\,
            I => \N__37338\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__37341\,
            I => acadc_skipcnt_15
        );

    \I__7112\ : Odrv4
    port map (
            O => \N__37338\,
            I => acadc_skipcnt_15
        );

    \I__7111\ : InMux
    port map (
            O => \N__37333\,
            I => \N__37330\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__37330\,
            I => \N__37326\
        );

    \I__7109\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37323\
        );

    \I__7108\ : Span4Mux_h
    port map (
            O => \N__37326\,
            I => \N__37320\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__37323\,
            I => acadc_skipcnt_9
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__37320\,
            I => acadc_skipcnt_9
        );

    \I__7105\ : InMux
    port map (
            O => \N__37315\,
            I => \N__37311\
        );

    \I__7104\ : InMux
    port map (
            O => \N__37314\,
            I => \N__37308\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__37311\,
            I => \N__37305\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__37308\,
            I => acadc_skipcnt_14
        );

    \I__7101\ : Odrv4
    port map (
            O => \N__37305\,
            I => acadc_skipcnt_14
        );

    \I__7100\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37296\
        );

    \I__7099\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37293\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__37296\,
            I => \N__37290\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__37293\,
            I => acadc_skipcnt_11
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__37290\,
            I => acadc_skipcnt_11
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__37285\,
            I => \N__37281\
        );

    \I__7094\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37276\
        );

    \I__7093\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37276\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__37276\,
            I => \N__37273\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__37273\,
            I => \N__37270\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__37270\,
            I => \N__37266\
        );

    \I__7089\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37263\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__37266\,
            I => cmd_rdadctmp_19
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__37263\,
            I => cmd_rdadctmp_19
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__37258\,
            I => \N__37255\
        );

    \I__7085\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37251\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__37254\,
            I => \N__37248\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37245\
        );

    \I__7082\ : InMux
    port map (
            O => \N__37248\,
            I => \N__37241\
        );

    \I__7081\ : Span4Mux_h
    port map (
            O => \N__37245\,
            I => \N__37238\
        );

    \I__7080\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37235\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__37241\,
            I => cmd_rdadctmp_20
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__37238\,
            I => cmd_rdadctmp_20
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__37235\,
            I => cmd_rdadctmp_20
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__37228\,
            I => \N__37224\
        );

    \I__7075\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37221\
        );

    \I__7074\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37217\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37214\
        );

    \I__7072\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37211\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37208\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__37214\,
            I => \N__37205\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__37211\,
            I => buf_dds1_0
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__37208\,
            I => buf_dds1_0
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__37205\,
            I => buf_dds1_0
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__37198\,
            I => \N__37195\
        );

    \I__7065\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37192\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37189\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__37189\,
            I => \N__37184\
        );

    \I__7062\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37181\
        );

    \I__7061\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37178\
        );

    \I__7060\ : Odrv4
    port map (
            O => \N__37184\,
            I => cmd_rdadctmp_28
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__37181\,
            I => cmd_rdadctmp_28
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__37178\,
            I => cmd_rdadctmp_28
        );

    \I__7057\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37168\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__37168\,
            I => \N__37165\
        );

    \I__7055\ : Span12Mux_s10_v
    port map (
            O => \N__37165\,
            I => \N__37160\
        );

    \I__7054\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37157\
        );

    \I__7053\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37154\
        );

    \I__7052\ : Span12Mux_v
    port map (
            O => \N__37160\,
            I => \N__37151\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37148\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__37154\,
            I => buf_adcdata_iac_20
        );

    \I__7049\ : Odrv12
    port map (
            O => \N__37151\,
            I => buf_adcdata_iac_20
        );

    \I__7048\ : Odrv4
    port map (
            O => \N__37148\,
            I => buf_adcdata_iac_20
        );

    \I__7047\ : SRMux
    port map (
            O => \N__37141\,
            I => \N__37138\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__37138\,
            I => \N__37135\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__37135\,
            I => \N__37131\
        );

    \I__7044\ : SRMux
    port map (
            O => \N__37134\,
            I => \N__37127\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__37131\,
            I => \N__37123\
        );

    \I__7042\ : SRMux
    port map (
            O => \N__37130\,
            I => \N__37120\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__37127\,
            I => \N__37117\
        );

    \I__7040\ : SRMux
    port map (
            O => \N__37126\,
            I => \N__37114\
        );

    \I__7039\ : Span4Mux_v
    port map (
            O => \N__37123\,
            I => \N__37109\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__37120\,
            I => \N__37109\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__37117\,
            I => \N__37104\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__37114\,
            I => \N__37104\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__37109\,
            I => \N__37101\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__37104\,
            I => \N__37098\
        );

    \I__7033\ : Span4Mux_v
    port map (
            O => \N__37101\,
            I => \N__37095\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__37098\,
            I => \N__37092\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__37095\,
            I => n15538
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__37092\,
            I => n15538
        );

    \I__7029\ : IoInMux
    port map (
            O => \N__37087\,
            I => \N__37084\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__37084\,
            I => \N__37080\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__37083\,
            I => \N__37076\
        );

    \I__7026\ : Span12Mux_s11_v
    port map (
            O => \N__37080\,
            I => \N__37073\
        );

    \I__7025\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37070\
        );

    \I__7024\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37067\
        );

    \I__7023\ : Odrv12
    port map (
            O => \N__37073\,
            I => \IAC_OSR0\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__37070\,
            I => \IAC_OSR0\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__37067\,
            I => \IAC_OSR0\
        );

    \I__7020\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__37057\,
            I => n24_adj_1575
        );

    \I__7018\ : IoInMux
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__7016\ : Span4Mux_s2_v
    port map (
            O => \N__37048\,
            I => \N__37044\
        );

    \I__7015\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37041\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__37044\,
            I => \N__37038\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__37041\,
            I => \N__37034\
        );

    \I__7012\ : Sp12to4
    port map (
            O => \N__37038\,
            I => \N__37031\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37028\
        );

    \I__7010\ : Span4Mux_h
    port map (
            O => \N__37034\,
            I => \N__37025\
        );

    \I__7009\ : Odrv12
    port map (
            O => \N__37031\,
            I => \IAC_OSR1\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__37028\,
            I => \IAC_OSR1\
        );

    \I__7007\ : Odrv4
    port map (
            O => \N__37025\,
            I => \IAC_OSR1\
        );

    \I__7006\ : InMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__37015\,
            I => n24_adj_1601
        );

    \I__7004\ : InMux
    port map (
            O => \N__37012\,
            I => \N__37009\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__37009\,
            I => n11984
        );

    \I__7002\ : InMux
    port map (
            O => \N__37006\,
            I => \N__37003\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__37003\,
            I => \N__37000\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__37000\,
            I => n16_adj_1733
        );

    \I__6999\ : InMux
    port map (
            O => \N__36997\,
            I => \N__36994\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__36994\,
            I => \N__36991\
        );

    \I__6997\ : Span12Mux_v
    port map (
            O => \N__36991\,
            I => \N__36988\
        );

    \I__6996\ : Odrv12
    port map (
            O => \N__36988\,
            I => n23438
        );

    \I__6995\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36982\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__36979\,
            I => \N__36974\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__36978\,
            I => \N__36971\
        );

    \I__6991\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36968\
        );

    \I__6990\ : Sp12to4
    port map (
            O => \N__36974\,
            I => \N__36965\
        );

    \I__6989\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36962\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__36968\,
            I => buf_adcdata_iac_12
        );

    \I__6987\ : Odrv12
    port map (
            O => \N__36965\,
            I => buf_adcdata_iac_12
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__36962\,
            I => buf_adcdata_iac_12
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__36955\,
            I => \N__36952\
        );

    \I__6984\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36948\
        );

    \I__6983\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36945\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__36948\,
            I => comm_test_buf_24_21
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__36945\,
            I => comm_test_buf_24_21
        );

    \I__6980\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36934\
        );

    \I__6978\ : Span4Mux_h
    port map (
            O => \N__36934\,
            I => \N__36930\
        );

    \I__6977\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36927\
        );

    \I__6976\ : Span4Mux_v
    port map (
            O => \N__36930\,
            I => \N__36922\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__36927\,
            I => \N__36922\
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__36922\,
            I => comm_test_buf_24_13
        );

    \I__6973\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36915\
        );

    \I__6972\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36911\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__36915\,
            I => \N__36908\
        );

    \I__6970\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36905\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__36911\,
            I => \N__36902\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__36908\,
            I => \N__36899\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36896\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__36902\,
            I => \N__36891\
        );

    \I__6965\ : Span4Mux_h
    port map (
            O => \N__36899\,
            I => \N__36891\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__36896\,
            I => \N__36888\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__36891\,
            I => comm_test_buf_24_5
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__36888\,
            I => comm_test_buf_24_5
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__36883\,
            I => \n111_adj_1776_cascade_\
        );

    \I__6960\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36877\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36874\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__36874\,
            I => \N__36871\
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__36871\,
            I => n111_adj_1761
        );

    \I__6956\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36864\
        );

    \I__6955\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36861\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__36864\,
            I => \N__36857\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__36861\,
            I => \N__36854\
        );

    \I__6952\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36851\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__36857\,
            I => \N__36846\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__36854\,
            I => \N__36846\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__36851\,
            I => buf_dds1_3
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__36846\,
            I => buf_dds1_3
        );

    \I__6947\ : InMux
    port map (
            O => \N__36841\,
            I => \N__36838\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__36838\,
            I => \N__36835\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__36835\,
            I => \N__36830\
        );

    \I__6944\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36825\
        );

    \I__6943\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36825\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__36830\,
            I => \N__36820\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__36825\,
            I => \N__36820\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__36820\,
            I => comm_buf_2_4
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__36817\,
            I => \n11987_cascade_\
        );

    \I__6938\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36811\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__36811\,
            I => \N__36808\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__36808\,
            I => \N__36805\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__36805\,
            I => n17_adj_1779
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__36802\,
            I => \n11985_cascade_\
        );

    \I__6933\ : CEMux
    port map (
            O => \N__36799\,
            I => \N__36795\
        );

    \I__6932\ : CEMux
    port map (
            O => \N__36798\,
            I => \N__36791\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__36795\,
            I => \N__36787\
        );

    \I__6930\ : CEMux
    port map (
            O => \N__36794\,
            I => \N__36784\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36781\
        );

    \I__6928\ : CEMux
    port map (
            O => \N__36790\,
            I => \N__36778\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__36787\,
            I => \N__36774\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36769\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__36781\,
            I => \N__36769\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__36778\,
            I => \N__36766\
        );

    \I__6923\ : InMux
    port map (
            O => \N__36777\,
            I => \N__36763\
        );

    \I__6922\ : Span4Mux_v
    port map (
            O => \N__36774\,
            I => \N__36760\
        );

    \I__6921\ : Span4Mux_v
    port map (
            O => \N__36769\,
            I => \N__36757\
        );

    \I__6920\ : Span4Mux_v
    port map (
            O => \N__36766\,
            I => \N__36752\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__36763\,
            I => \N__36752\
        );

    \I__6918\ : Span4Mux_v
    port map (
            O => \N__36760\,
            I => \N__36749\
        );

    \I__6917\ : Sp12to4
    port map (
            O => \N__36757\,
            I => \N__36746\
        );

    \I__6916\ : Span4Mux_v
    port map (
            O => \N__36752\,
            I => \N__36743\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__36749\,
            I => \N__36740\
        );

    \I__6914\ : Span12Mux_v
    port map (
            O => \N__36746\,
            I => \N__36737\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__36743\,
            I => \N__36734\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__36740\,
            I => n13117
        );

    \I__6911\ : Odrv12
    port map (
            O => \N__36737\,
            I => n13117
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__36734\,
            I => n13117
        );

    \I__6909\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36724\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__36724\,
            I => \N__36721\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__36721\,
            I => \N__36718\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__36718\,
            I => \comm_buf_2_7_N_575_7\
        );

    \I__6905\ : SRMux
    port map (
            O => \N__36715\,
            I => \N__36712\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__36712\,
            I => \N__36709\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__36709\,
            I => \N__36706\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__6901\ : Odrv4
    port map (
            O => \N__36703\,
            I => \comm_spi.data_tx_7__N_859\
        );

    \I__6900\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36675\
        );

    \I__6899\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36675\
        );

    \I__6898\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36675\
        );

    \I__6897\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36675\
        );

    \I__6896\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36675\
        );

    \I__6895\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36675\
        );

    \I__6894\ : InMux
    port map (
            O => \N__36694\,
            I => \N__36675\
        );

    \I__6893\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36675\
        );

    \I__6892\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36672\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__36675\,
            I => \N__36662\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36659\
        );

    \I__6889\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36644\
        );

    \I__6888\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36644\
        );

    \I__6887\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36644\
        );

    \I__6886\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36644\
        );

    \I__6885\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36644\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36644\
        );

    \I__6883\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36644\
        );

    \I__6882\ : Sp12to4
    port map (
            O => \N__36662\,
            I => \N__36641\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__36659\,
            I => n6774
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__36644\,
            I => n6774
        );

    \I__6879\ : Odrv12
    port map (
            O => \N__36641\,
            I => n6774
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__36634\,
            I => \n111_adj_1796_cascade_\
        );

    \I__6877\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36625\
        );

    \I__6876\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36625\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__36625\,
            I => comm_test_buf_24_10
        );

    \I__6874\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36619\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__36619\,
            I => \N__36616\
        );

    \I__6872\ : Span4Mux_v
    port map (
            O => \N__36616\,
            I => \N__36612\
        );

    \I__6871\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36609\
        );

    \I__6870\ : Span4Mux_h
    port map (
            O => \N__36612\,
            I => \N__36606\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36603\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__36606\,
            I => \comm_spi.n15365\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__36603\,
            I => \comm_spi.n15365\
        );

    \I__6866\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36595\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__36595\,
            I => \N__36592\
        );

    \I__6864\ : Span4Mux_v
    port map (
            O => \N__36592\,
            I => \N__36587\
        );

    \I__6863\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36584\
        );

    \I__6862\ : InMux
    port map (
            O => \N__36590\,
            I => \N__36581\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__36587\,
            I => \comm_spi.n24025\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__36584\,
            I => \comm_spi.n24025\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__36581\,
            I => \comm_spi.n24025\
        );

    \I__6858\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36571\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__36571\,
            I => \N__36568\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__36568\,
            I => \N__36565\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__36565\,
            I => \N__36561\
        );

    \I__6854\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36558\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__36561\,
            I => \comm_spi.n15364\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__36558\,
            I => \comm_spi.n15364\
        );

    \I__6851\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36549\
        );

    \I__6850\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36546\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36543\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__36546\,
            I => \N__36540\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__36543\,
            I => \N__36535\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__36540\,
            I => \N__36535\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__36535\,
            I => \N__36532\
        );

    \I__6844\ : Odrv4
    port map (
            O => \N__36532\,
            I => \comm_spi.n15368\
        );

    \I__6843\ : SRMux
    port map (
            O => \N__36529\,
            I => \N__36526\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__36526\,
            I => \N__36523\
        );

    \I__6841\ : Span4Mux_v
    port map (
            O => \N__36523\,
            I => \N__36520\
        );

    \I__6840\ : Span4Mux_v
    port map (
            O => \N__36520\,
            I => \N__36517\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__36517\,
            I => \comm_spi.data_tx_7__N_855\
        );

    \I__6838\ : IoInMux
    port map (
            O => \N__36514\,
            I => \N__36511\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36508\
        );

    \I__6836\ : Span4Mux_s2_h
    port map (
            O => \N__36508\,
            I => \N__36505\
        );

    \I__6835\ : Span4Mux_v
    port map (
            O => \N__36505\,
            I => \N__36502\
        );

    \I__6834\ : Sp12to4
    port map (
            O => \N__36502\,
            I => \N__36497\
        );

    \I__6833\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36494\
        );

    \I__6832\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36491\
        );

    \I__6831\ : Span12Mux_h
    port map (
            O => \N__36497\,
            I => \N__36486\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__36494\,
            I => \N__36486\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__36491\,
            I => \AMPV_POW\
        );

    \I__6828\ : Odrv12
    port map (
            O => \N__36486\,
            I => \AMPV_POW\
        );

    \I__6827\ : CascadeMux
    port map (
            O => \N__36481\,
            I => \N__36478\
        );

    \I__6826\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36475\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__36475\,
            I => \N__36472\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__36472\,
            I => \N__36469\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__36469\,
            I => \comm_buf_0_7_N_543_7\
        );

    \I__6822\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36462\
        );

    \I__6821\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36459\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__36462\,
            I => \N__36455\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__36459\,
            I => \N__36452\
        );

    \I__6818\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36449\
        );

    \I__6817\ : Span4Mux_v
    port map (
            O => \N__36455\,
            I => \N__36446\
        );

    \I__6816\ : Odrv4
    port map (
            O => \N__36452\,
            I => clk_cnt_1
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__36449\,
            I => clk_cnt_1
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__36446\,
            I => clk_cnt_1
        );

    \I__6813\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36433\
        );

    \I__6812\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36430\
        );

    \I__6811\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36425\
        );

    \I__6810\ : InMux
    port map (
            O => \N__36436\,
            I => \N__36425\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__36433\,
            I => \N__36420\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__36430\,
            I => \N__36420\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__36425\,
            I => clk_cnt_0
        );

    \I__6806\ : Odrv12
    port map (
            O => \N__36420\,
            I => clk_cnt_0
        );

    \I__6805\ : SRMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36409\
        );

    \I__6803\ : Span4Mux_v
    port map (
            O => \N__36409\,
            I => \N__36406\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__36406\,
            I => \N__36403\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__36403\,
            I => n18996
        );

    \I__6800\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36397\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__36397\,
            I => \comm_buf_2_7_N_575_0\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__36394\,
            I => \N__36391\
        );

    \I__6797\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36388\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36385\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__36385\,
            I => \comm_buf_2_7_N_575_1\
        );

    \I__6794\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36379\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__36379\,
            I => \N__36376\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__36376\,
            I => \comm_buf_2_7_N_575_3\
        );

    \I__6791\ : InMux
    port map (
            O => \N__36373\,
            I => \N__36370\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__36370\,
            I => \N__36367\
        );

    \I__6789\ : Odrv12
    port map (
            O => \N__36367\,
            I => \comm_buf_2_7_N_575_4\
        );

    \I__6788\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36361\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__36361\,
            I => \N__36358\
        );

    \I__6786\ : Odrv12
    port map (
            O => \N__36358\,
            I => \comm_buf_2_7_N_575_5\
        );

    \I__6785\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36352\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36349\
        );

    \I__6783\ : Odrv12
    port map (
            O => \N__36349\,
            I => \comm_buf_2_7_N_575_6\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__36346\,
            I => \N__36343\
        );

    \I__6781\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36338\
        );

    \I__6780\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36333\
        );

    \I__6779\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36333\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__36338\,
            I => \N__36330\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__36333\,
            I => \N__36327\
        );

    \I__6776\ : Span4Mux_h
    port map (
            O => \N__36330\,
            I => \N__36324\
        );

    \I__6775\ : Sp12to4
    port map (
            O => \N__36327\,
            I => \N__36321\
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__36324\,
            I => comm_buf_2_6
        );

    \I__6773\ : Odrv12
    port map (
            O => \N__36321\,
            I => comm_buf_2_6
        );

    \I__6772\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36313\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__36313\,
            I => n22669
        );

    \I__6770\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36307\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__36304\,
            I => n1_adj_1668
        );

    \I__6767\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36298\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__36298\,
            I => n13219
        );

    \I__6765\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36289\
        );

    \I__6764\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36289\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__36289\,
            I => \N__36286\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__36286\,
            I => \N__36282\
        );

    \I__6761\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36279\
        );

    \I__6760\ : Odrv4
    port map (
            O => \N__36282\,
            I => comm_tx_buf_4
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__36279\,
            I => comm_tx_buf_4
        );

    \I__6758\ : SRMux
    port map (
            O => \N__36274\,
            I => \N__36271\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__36268\,
            I => \N__36265\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__36265\,
            I => \comm_spi.data_tx_7__N_871\
        );

    \I__6754\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36259\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__36259\,
            I => \N__36256\
        );

    \I__6752\ : Odrv12
    port map (
            O => \N__36256\,
            I => \comm_buf_0_7_N_543_4\
        );

    \I__6751\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36250\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N__36247\
        );

    \I__6749\ : Span4Mux_h
    port map (
            O => \N__36247\,
            I => \N__36244\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__36244\,
            I => \comm_buf_0_7_N_543_6\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__36241\,
            I => \comm_spi.n24034_cascade_\
        );

    \I__6746\ : InMux
    port map (
            O => \N__36238\,
            I => \N__36235\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__36235\,
            I => \N__36232\
        );

    \I__6744\ : Span4Mux_h
    port map (
            O => \N__36232\,
            I => \N__36228\
        );

    \I__6743\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36225\
        );

    \I__6742\ : Span4Mux_h
    port map (
            O => \N__36228\,
            I => \N__36222\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36219\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__36222\,
            I => \comm_spi.n15356\
        );

    \I__6739\ : Odrv4
    port map (
            O => \N__36219\,
            I => \comm_spi.n15356\
        );

    \I__6738\ : SRMux
    port map (
            O => \N__36214\,
            I => \N__36211\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__36211\,
            I => \N__36208\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__36208\,
            I => \N__36205\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__36205\,
            I => \comm_spi.data_tx_7__N_858\
        );

    \I__6734\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36195\
        );

    \I__6733\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36195\
        );

    \I__6732\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36192\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36195\,
            I => comm_tx_buf_6
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__36192\,
            I => comm_tx_buf_6
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__36187\,
            I => \N__36184\
        );

    \I__6728\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36180\
        );

    \I__6727\ : InMux
    port map (
            O => \N__36183\,
            I => \N__36177\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__36180\,
            I => \N__36172\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36172\
        );

    \I__6724\ : Span4Mux_v
    port map (
            O => \N__36172\,
            I => \N__36169\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__36169\,
            I => \N__36165\
        );

    \I__6722\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36162\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__36165\,
            I => \comm_spi.n24013\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__36162\,
            I => \comm_spi.n24013\
        );

    \I__6719\ : SRMux
    port map (
            O => \N__36157\,
            I => \N__36154\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__36154\,
            I => \N__36151\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__36151\,
            I => \N__36148\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__36148\,
            I => \N__36145\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__36145\,
            I => \comm_spi.data_tx_7__N_856\
        );

    \I__6714\ : CascadeMux
    port map (
            O => \N__36142\,
            I => \n2_adj_1669_cascade_\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__36139\,
            I => \n4_adj_1670_cascade_\
        );

    \I__6712\ : InMux
    port map (
            O => \N__36136\,
            I => \N__36133\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__36133\,
            I => n23402
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__36130\,
            I => \n19_adj_1706_cascade_\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__36127\,
            I => \N__36123\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__36126\,
            I => \N__36120\
        );

    \I__6707\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36117\
        );

    \I__6706\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36114\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__36110\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36107\
        );

    \I__6703\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36104\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__36110\,
            I => \N__36101\
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__36107\,
            I => cmd_rdadctmp_8_adj_1540
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__36104\,
            I => cmd_rdadctmp_8_adj_1540
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__36101\,
            I => cmd_rdadctmp_8_adj_1540
        );

    \I__6698\ : InMux
    port map (
            O => \N__36094\,
            I => \N__36090\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__36093\,
            I => \N__36087\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36083\
        );

    \I__6695\ : InMux
    port map (
            O => \N__36087\,
            I => \N__36080\
        );

    \I__6694\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36077\
        );

    \I__6693\ : Span12Mux_h
    port map (
            O => \N__36083\,
            I => \N__36074\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__36080\,
            I => buf_adcdata_iac_1
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__36077\,
            I => buf_adcdata_iac_1
        );

    \I__6690\ : Odrv12
    port map (
            O => \N__36074\,
            I => buf_adcdata_iac_1
        );

    \I__6689\ : InMux
    port map (
            O => \N__36067\,
            I => \N__36064\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__36061\
        );

    \I__6687\ : Span4Mux_v
    port map (
            O => \N__36061\,
            I => \N__36058\
        );

    \I__6686\ : Sp12to4
    port map (
            O => \N__36058\,
            I => \N__36053\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36048\
        );

    \I__6684\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36048\
        );

    \I__6683\ : Odrv12
    port map (
            O => \N__36053\,
            I => buf_adcdata_iac_2
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__36048\,
            I => buf_adcdata_iac_2
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__36043\,
            I => \N__36040\
        );

    \I__6680\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36037\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__36037\,
            I => \N__36034\
        );

    \I__6678\ : Span4Mux_h
    port map (
            O => \N__36034\,
            I => \N__36030\
        );

    \I__6677\ : InMux
    port map (
            O => \N__36033\,
            I => \N__36026\
        );

    \I__6676\ : Span4Mux_h
    port map (
            O => \N__36030\,
            I => \N__36023\
        );

    \I__6675\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36020\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__36026\,
            I => cmd_rdadctmp_10_adj_1538
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__36023\,
            I => cmd_rdadctmp_10_adj_1538
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__36020\,
            I => cmd_rdadctmp_10_adj_1538
        );

    \I__6671\ : InMux
    port map (
            O => \N__36013\,
            I => \N__35994\
        );

    \I__6670\ : InMux
    port map (
            O => \N__36012\,
            I => \N__35977\
        );

    \I__6669\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35977\
        );

    \I__6668\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35977\
        );

    \I__6667\ : InMux
    port map (
            O => \N__36009\,
            I => \N__35977\
        );

    \I__6666\ : InMux
    port map (
            O => \N__36008\,
            I => \N__35977\
        );

    \I__6665\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35966\
        );

    \I__6664\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35966\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35966\
        );

    \I__6662\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35966\
        );

    \I__6661\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35966\
        );

    \I__6660\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35959\
        );

    \I__6659\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35947\
        );

    \I__6658\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35947\
        );

    \I__6657\ : InMux
    port map (
            O => \N__35999\,
            I => \N__35947\
        );

    \I__6656\ : InMux
    port map (
            O => \N__35998\,
            I => \N__35947\
        );

    \I__6655\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35947\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__35994\,
            I => \N__35943\
        );

    \I__6653\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35938\
        );

    \I__6652\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35938\
        );

    \I__6651\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35933\
        );

    \I__6650\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35933\
        );

    \I__6649\ : CascadeMux
    port map (
            O => \N__35989\,
            I => \N__35930\
        );

    \I__6648\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35918\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__35977\,
            I => \N__35904\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__35966\,
            I => \N__35904\
        );

    \I__6645\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35899\
        );

    \I__6644\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35899\
        );

    \I__6643\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35891\
        );

    \I__6642\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35891\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35888\
        );

    \I__6640\ : InMux
    port map (
            O => \N__35958\,
            I => \N__35885\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__35947\,
            I => \N__35882\
        );

    \I__6638\ : InMux
    port map (
            O => \N__35946\,
            I => \N__35878\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__35943\,
            I => \N__35875\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35872\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35869\
        );

    \I__6634\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35860\
        );

    \I__6633\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35860\
        );

    \I__6632\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35855\
        );

    \I__6631\ : InMux
    port map (
            O => \N__35927\,
            I => \N__35855\
        );

    \I__6630\ : InMux
    port map (
            O => \N__35926\,
            I => \N__35851\
        );

    \I__6629\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35846\
        );

    \I__6628\ : InMux
    port map (
            O => \N__35924\,
            I => \N__35846\
        );

    \I__6627\ : InMux
    port map (
            O => \N__35923\,
            I => \N__35843\
        );

    \I__6626\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35838\
        );

    \I__6625\ : InMux
    port map (
            O => \N__35921\,
            I => \N__35838\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__35918\,
            I => \N__35835\
        );

    \I__6623\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35826\
        );

    \I__6622\ : InMux
    port map (
            O => \N__35916\,
            I => \N__35826\
        );

    \I__6621\ : InMux
    port map (
            O => \N__35915\,
            I => \N__35826\
        );

    \I__6620\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35826\
        );

    \I__6619\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35819\
        );

    \I__6618\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35819\
        );

    \I__6617\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35819\
        );

    \I__6616\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35814\
        );

    \I__6615\ : InMux
    port map (
            O => \N__35909\,
            I => \N__35814\
        );

    \I__6614\ : Span4Mux_v
    port map (
            O => \N__35904\,
            I => \N__35809\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35809\
        );

    \I__6612\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35802\
        );

    \I__6611\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35802\
        );

    \I__6610\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35802\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35799\
        );

    \I__6608\ : Span4Mux_v
    port map (
            O => \N__35888\,
            I => \N__35792\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__35885\,
            I => \N__35792\
        );

    \I__6606\ : Span4Mux_h
    port map (
            O => \N__35882\,
            I => \N__35792\
        );

    \I__6605\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35789\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35786\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__35875\,
            I => \N__35779\
        );

    \I__6602\ : Span4Mux_v
    port map (
            O => \N__35872\,
            I => \N__35779\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__35869\,
            I => \N__35779\
        );

    \I__6600\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35771\
        );

    \I__6599\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35768\
        );

    \I__6598\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35763\
        );

    \I__6597\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35763\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__35860\,
            I => \N__35758\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35758\
        );

    \I__6594\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35755\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__35851\,
            I => \N__35748\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35748\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35748\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35745\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__35835\,
            I => \N__35740\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__35826\,
            I => \N__35740\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__35819\,
            I => \N__35737\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35730\
        );

    \I__6585\ : Span4Mux_h
    port map (
            O => \N__35809\,
            I => \N__35730\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__35802\,
            I => \N__35730\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__35799\,
            I => \N__35727\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__35792\,
            I => \N__35724\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35717\
        );

    \I__6580\ : Span4Mux_h
    port map (
            O => \N__35786\,
            I => \N__35717\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__35779\,
            I => \N__35717\
        );

    \I__6578\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35702\
        );

    \I__6577\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35702\
        );

    \I__6576\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35702\
        );

    \I__6575\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35697\
        );

    \I__6574\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35697\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35692\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35692\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__35763\,
            I => \N__35687\
        );

    \I__6570\ : Span12Mux_h
    port map (
            O => \N__35758\,
            I => \N__35687\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35670\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35670\
        );

    \I__6567\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35670\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__35740\,
            I => \N__35670\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__35737\,
            I => \N__35670\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__35730\,
            I => \N__35670\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__35727\,
            I => \N__35670\
        );

    \I__6562\ : Span4Mux_h
    port map (
            O => \N__35724\,
            I => \N__35670\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__35717\,
            I => \N__35667\
        );

    \I__6560\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35662\
        );

    \I__6559\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35662\
        );

    \I__6558\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35653\
        );

    \I__6557\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35653\
        );

    \I__6556\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35653\
        );

    \I__6555\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35653\
        );

    \I__6554\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35648\
        );

    \I__6553\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35648\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__35702\,
            I => adc_state_0_adj_1516
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__35697\,
            I => adc_state_0_adj_1516
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__35692\,
            I => adc_state_0_adj_1516
        );

    \I__6549\ : Odrv12
    port map (
            O => \N__35687\,
            I => adc_state_0_adj_1516
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__35670\,
            I => adc_state_0_adj_1516
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__35667\,
            I => adc_state_0_adj_1516
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__35662\,
            I => adc_state_0_adj_1516
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__35653\,
            I => adc_state_0_adj_1516
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__35648\,
            I => adc_state_0_adj_1516
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__35629\,
            I => \N__35626\
        );

    \I__6542\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35618\
        );

    \I__6541\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35618\
        );

    \I__6540\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35611\
        );

    \I__6539\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35611\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__35618\,
            I => \N__35604\
        );

    \I__6537\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35591\
        );

    \I__6536\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35591\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__35611\,
            I => \N__35588\
        );

    \I__6534\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35584\
        );

    \I__6533\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35581\
        );

    \I__6532\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35578\
        );

    \I__6531\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35575\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__35604\,
            I => \N__35572\
        );

    \I__6529\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35568\
        );

    \I__6528\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35562\
        );

    \I__6527\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35559\
        );

    \I__6526\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35552\
        );

    \I__6525\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35552\
        );

    \I__6524\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35552\
        );

    \I__6523\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35547\
        );

    \I__6522\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35547\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35542\
        );

    \I__6520\ : Span4Mux_v
    port map (
            O => \N__35588\,
            I => \N__35542\
        );

    \I__6519\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35539\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35534\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__35581\,
            I => \N__35534\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__35578\,
            I => \N__35531\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__35575\,
            I => \N__35526\
        );

    \I__6514\ : Span4Mux_h
    port map (
            O => \N__35572\,
            I => \N__35526\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35523\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35520\
        );

    \I__6511\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35517\
        );

    \I__6510\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35512\
        );

    \I__6509\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35512\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35507\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35507\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__35552\,
            I => \N__35504\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35499\
        );

    \I__6504\ : Span4Mux_h
    port map (
            O => \N__35542\,
            I => \N__35499\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35494\
        );

    \I__6502\ : Span4Mux_v
    port map (
            O => \N__35534\,
            I => \N__35494\
        );

    \I__6501\ : Span4Mux_v
    port map (
            O => \N__35531\,
            I => \N__35489\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__35526\,
            I => \N__35489\
        );

    \I__6499\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35486\
        );

    \I__6498\ : Span4Mux_h
    port map (
            O => \N__35520\,
            I => \N__35483\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__35517\,
            I => \N__35472\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35472\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__35507\,
            I => \N__35472\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__35504\,
            I => \N__35472\
        );

    \I__6493\ : Span4Mux_h
    port map (
            O => \N__35499\,
            I => \N__35472\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__35494\,
            I => \N__35467\
        );

    \I__6491\ : Span4Mux_h
    port map (
            O => \N__35489\,
            I => \N__35467\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__35486\,
            I => n21948
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__35483\,
            I => n21948
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__35472\,
            I => n21948
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__35467\,
            I => n21948
        );

    \I__6486\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35455\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__35455\,
            I => \N__35452\
        );

    \I__6484\ : Span4Mux_v
    port map (
            O => \N__35452\,
            I => \N__35449\
        );

    \I__6483\ : Sp12to4
    port map (
            O => \N__35449\,
            I => \N__35444\
        );

    \I__6482\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35439\
        );

    \I__6481\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35439\
        );

    \I__6480\ : Odrv12
    port map (
            O => \N__35444\,
            I => buf_adcdata_vac_2
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__35439\,
            I => buf_adcdata_vac_2
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__35434\,
            I => \N__35430\
        );

    \I__6477\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35425\
        );

    \I__6476\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35425\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__35425\,
            I => \N__35422\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__35422\,
            I => \N__35418\
        );

    \I__6473\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35415\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__35418\,
            I => cmd_rdadctmp_9
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__35415\,
            I => cmd_rdadctmp_9
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__35410\,
            I => \N__35406\
        );

    \I__6469\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35398\
        );

    \I__6468\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35398\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35398\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__35398\,
            I => cmd_rdadctmp_10
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__35395\,
            I => \N__35392\
        );

    \I__6464\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35389\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__35389\,
            I => \N__35385\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__35388\,
            I => \N__35382\
        );

    \I__6461\ : Span4Mux_v
    port map (
            O => \N__35385\,
            I => \N__35379\
        );

    \I__6460\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35375\
        );

    \I__6459\ : Span4Mux_h
    port map (
            O => \N__35379\,
            I => \N__35372\
        );

    \I__6458\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35369\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__35375\,
            I => cmd_rdadctmp_11
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__35372\,
            I => cmd_rdadctmp_11
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__35369\,
            I => cmd_rdadctmp_11
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__35362\,
            I => \N__35359\
        );

    \I__6453\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35356\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__35356\,
            I => \N__35351\
        );

    \I__6451\ : InMux
    port map (
            O => \N__35355\,
            I => \N__35348\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__35354\,
            I => \N__35345\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__35351\,
            I => \N__35341\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__35348\,
            I => \N__35338\
        );

    \I__6447\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35334\
        );

    \I__6446\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35331\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__35341\,
            I => \N__35326\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__35338\,
            I => \N__35326\
        );

    \I__6443\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35323\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35318\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__35331\,
            I => \N__35318\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__35326\,
            I => \buf_cfgRTD_7\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__35323\,
            I => \buf_cfgRTD_7\
        );

    \I__6438\ : Odrv12
    port map (
            O => \N__35318\,
            I => \buf_cfgRTD_7\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__35311\,
            I => \N__35308\
        );

    \I__6436\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35305\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__35305\,
            I => \N__35302\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__35302\,
            I => \N__35299\
        );

    \I__6433\ : Span4Mux_h
    port map (
            O => \N__35299\,
            I => \N__35295\
        );

    \I__6432\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35292\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__35295\,
            I => \buf_readRTD_15\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__35292\,
            I => \buf_readRTD_15\
        );

    \I__6429\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35284\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__35284\,
            I => \N__35281\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__35281\,
            I => \N__35278\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__35278\,
            I => n23432
        );

    \I__6425\ : CascadeMux
    port map (
            O => \N__35275\,
            I => \n12610_cascade_\
        );

    \I__6424\ : SRMux
    port map (
            O => \N__35272\,
            I => \N__35269\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__35269\,
            I => \N__35266\
        );

    \I__6422\ : Span4Mux_h
    port map (
            O => \N__35266\,
            I => \N__35263\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__35263\,
            I => \N__35260\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__35260\,
            I => \comm_spi.data_tx_7__N_883\
        );

    \I__6419\ : IoInMux
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35251\
        );

    \I__6417\ : Span4Mux_s3_h
    port map (
            O => \N__35251\,
            I => \N__35248\
        );

    \I__6416\ : Span4Mux_v
    port map (
            O => \N__35248\,
            I => \N__35245\
        );

    \I__6415\ : Sp12to4
    port map (
            O => \N__35245\,
            I => \N__35242\
        );

    \I__6414\ : Span12Mux_h
    port map (
            O => \N__35242\,
            I => \N__35239\
        );

    \I__6413\ : Odrv12
    port map (
            O => \N__35239\,
            I => \ICE_SPI_MISO\
        );

    \I__6412\ : SRMux
    port map (
            O => \N__35236\,
            I => \N__35233\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__35233\,
            I => \N__35230\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__35224\,
            I => \comm_spi.data_tx_7__N_868\
        );

    \I__6407\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35218\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__6405\ : Span4Mux_h
    port map (
            O => \N__35215\,
            I => \N__35211\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__35214\,
            I => \N__35208\
        );

    \I__6403\ : Span4Mux_v
    port map (
            O => \N__35211\,
            I => \N__35205\
        );

    \I__6402\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35202\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__35205\,
            I => buf_adcdata_vdc_2
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__35202\,
            I => buf_adcdata_vdc_2
        );

    \I__6399\ : InMux
    port map (
            O => \N__35197\,
            I => n20649
        );

    \I__6398\ : InMux
    port map (
            O => \N__35194\,
            I => n20650
        );

    \I__6397\ : InMux
    port map (
            O => \N__35191\,
            I => n20651
        );

    \I__6396\ : CEMux
    port map (
            O => \N__35188\,
            I => \N__35184\
        );

    \I__6395\ : CEMux
    port map (
            O => \N__35187\,
            I => \N__35181\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__35184\,
            I => \N__35178\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__35181\,
            I => \N__35175\
        );

    \I__6392\ : Span4Mux_v
    port map (
            O => \N__35178\,
            I => \N__35172\
        );

    \I__6391\ : Span4Mux_v
    port map (
            O => \N__35175\,
            I => \N__35168\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__35172\,
            I => \N__35165\
        );

    \I__6389\ : CEMux
    port map (
            O => \N__35171\,
            I => \N__35162\
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__35168\,
            I => n12450
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__35165\,
            I => n12450
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__35162\,
            I => n12450
        );

    \I__6385\ : SRMux
    port map (
            O => \N__35155\,
            I => \N__35151\
        );

    \I__6384\ : SRMux
    port map (
            O => \N__35154\,
            I => \N__35148\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35145\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__35148\,
            I => \N__35142\
        );

    \I__6381\ : Span4Mux_v
    port map (
            O => \N__35145\,
            I => \N__35139\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__35142\,
            I => \N__35136\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__35139\,
            I => n15439
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__35136\,
            I => n15439
        );

    \I__6377\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35125\
        );

    \I__6376\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35118\
        );

    \I__6375\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35118\
        );

    \I__6374\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35118\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35112\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__35112\
        );

    \I__6371\ : InMux
    port map (
            O => \N__35117\,
            I => \N__35109\
        );

    \I__6370\ : Span12Mux_s11_h
    port map (
            O => \N__35112\,
            I => \N__35106\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__35109\,
            I => \RTD.bit_cnt_3\
        );

    \I__6368\ : Odrv12
    port map (
            O => \N__35106\,
            I => \RTD.bit_cnt_3\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__35101\,
            I => \N__35098\
        );

    \I__6366\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35091\
        );

    \I__6365\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35091\
        );

    \I__6364\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35088\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__35091\,
            I => \RTD.bit_cnt_2\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__35088\,
            I => \RTD.bit_cnt_2\
        );

    \I__6361\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35073\
        );

    \I__6360\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35073\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35073\
        );

    \I__6358\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35070\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__35073\,
            I => \RTD.bit_cnt_1\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__35070\,
            I => \RTD.bit_cnt_1\
        );

    \I__6355\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35052\
        );

    \I__6354\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35052\
        );

    \I__6353\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35052\
        );

    \I__6352\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35052\
        );

    \I__6351\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35049\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__35052\,
            I => \RTD.bit_cnt_0\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__35049\,
            I => \RTD.bit_cnt_0\
        );

    \I__6348\ : ClkMux
    port map (
            O => \N__35044\,
            I => \N__35039\
        );

    \I__6347\ : ClkMux
    port map (
            O => \N__35043\,
            I => \N__35035\
        );

    \I__6346\ : ClkMux
    port map (
            O => \N__35042\,
            I => \N__35031\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__35039\,
            I => \N__35026\
        );

    \I__6344\ : ClkMux
    port map (
            O => \N__35038\,
            I => \N__35023\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35018\
        );

    \I__6342\ : ClkMux
    port map (
            O => \N__35034\,
            I => \N__35015\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35010\
        );

    \I__6340\ : ClkMux
    port map (
            O => \N__35030\,
            I => \N__35007\
        );

    \I__6339\ : ClkMux
    port map (
            O => \N__35029\,
            I => \N__35003\
        );

    \I__6338\ : Span4Mux_h
    port map (
            O => \N__35026\,
            I => \N__34995\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__34995\
        );

    \I__6336\ : ClkMux
    port map (
            O => \N__35022\,
            I => \N__34992\
        );

    \I__6335\ : ClkMux
    port map (
            O => \N__35021\,
            I => \N__34989\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__35018\,
            I => \N__34984\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__34984\
        );

    \I__6332\ : ClkMux
    port map (
            O => \N__35014\,
            I => \N__34981\
        );

    \I__6331\ : ClkMux
    port map (
            O => \N__35013\,
            I => \N__34977\
        );

    \I__6330\ : Span4Mux_h
    port map (
            O => \N__35010\,
            I => \N__34972\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__35007\,
            I => \N__34972\
        );

    \I__6328\ : ClkMux
    port map (
            O => \N__35006\,
            I => \N__34969\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__35003\,
            I => \N__34966\
        );

    \I__6326\ : ClkMux
    port map (
            O => \N__35002\,
            I => \N__34963\
        );

    \I__6325\ : ClkMux
    port map (
            O => \N__35001\,
            I => \N__34960\
        );

    \I__6324\ : ClkMux
    port map (
            O => \N__35000\,
            I => \N__34957\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__34995\,
            I => \N__34953\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__34992\,
            I => \N__34948\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__34989\,
            I => \N__34948\
        );

    \I__6320\ : Span4Mux_v
    port map (
            O => \N__34984\,
            I => \N__34943\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__34981\,
            I => \N__34943\
        );

    \I__6318\ : ClkMux
    port map (
            O => \N__34980\,
            I => \N__34940\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__34977\,
            I => \N__34937\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__34972\,
            I => \N__34932\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34932\
        );

    \I__6314\ : Span4Mux_h
    port map (
            O => \N__34966\,
            I => \N__34927\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34927\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34924\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__34957\,
            I => \N__34921\
        );

    \I__6310\ : ClkMux
    port map (
            O => \N__34956\,
            I => \N__34918\
        );

    \I__6309\ : Span4Mux_h
    port map (
            O => \N__34953\,
            I => \N__34909\
        );

    \I__6308\ : Span4Mux_v
    port map (
            O => \N__34948\,
            I => \N__34909\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__34943\,
            I => \N__34909\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34909\
        );

    \I__6305\ : Span4Mux_v
    port map (
            O => \N__34937\,
            I => \N__34902\
        );

    \I__6304\ : Span4Mux_h
    port map (
            O => \N__34932\,
            I => \N__34902\
        );

    \I__6303\ : Span4Mux_v
    port map (
            O => \N__34927\,
            I => \N__34902\
        );

    \I__6302\ : Span4Mux_v
    port map (
            O => \N__34924\,
            I => \N__34895\
        );

    \I__6301\ : Span4Mux_v
    port map (
            O => \N__34921\,
            I => \N__34895\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34895\
        );

    \I__6299\ : Span4Mux_h
    port map (
            O => \N__34909\,
            I => \N__34892\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__34902\,
            I => \N__34887\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__34895\,
            I => \N__34887\
        );

    \I__6296\ : Span4Mux_h
    port map (
            O => \N__34892\,
            I => \N__34882\
        );

    \I__6295\ : Span4Mux_h
    port map (
            O => \N__34887\,
            I => \N__34879\
        );

    \I__6294\ : ClkMux
    port map (
            O => \N__34886\,
            I => \N__34876\
        );

    \I__6293\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34873\
        );

    \I__6292\ : Odrv4
    port map (
            O => \N__34882\,
            I => \clk_RTD\
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__34879\,
            I => \clk_RTD\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__34876\,
            I => \clk_RTD\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__34873\,
            I => \clk_RTD\
        );

    \I__6288\ : CEMux
    port map (
            O => \N__34864\,
            I => \N__34861\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34858\
        );

    \I__6286\ : Span4Mux_h
    port map (
            O => \N__34858\,
            I => \N__34855\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__34855\,
            I => \RTD.n18274\
        );

    \I__6284\ : SRMux
    port map (
            O => \N__34852\,
            I => \N__34849\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__34849\,
            I => \N__34846\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__34846\,
            I => \N__34843\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__34843\,
            I => \RTD.n18275\
        );

    \I__6280\ : InMux
    port map (
            O => \N__34840\,
            I => n20640
        );

    \I__6279\ : InMux
    port map (
            O => \N__34837\,
            I => n20641
        );

    \I__6278\ : InMux
    port map (
            O => \N__34834\,
            I => n20642
        );

    \I__6277\ : InMux
    port map (
            O => \N__34831\,
            I => n20643
        );

    \I__6276\ : InMux
    port map (
            O => \N__34828\,
            I => n20644
        );

    \I__6275\ : InMux
    port map (
            O => \N__34825\,
            I => \bfn_11_20_0_\
        );

    \I__6274\ : InMux
    port map (
            O => \N__34822\,
            I => n20646
        );

    \I__6273\ : InMux
    port map (
            O => \N__34819\,
            I => n20647
        );

    \I__6272\ : InMux
    port map (
            O => \N__34816\,
            I => n20648
        );

    \I__6271\ : InMux
    port map (
            O => \N__34813\,
            I => \bfn_11_19_0_\
        );

    \I__6270\ : InMux
    port map (
            O => \N__34810\,
            I => n20638
        );

    \I__6269\ : InMux
    port map (
            O => \N__34807\,
            I => n20639
        );

    \I__6268\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34801\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__34801\,
            I => n11980
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__34798\,
            I => \N__34792\
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__34797\,
            I => \N__34788\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__34796\,
            I => \N__34778\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34775\
        );

    \I__6262\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34771\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__34791\,
            I => \N__34768\
        );

    \I__6260\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34765\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__34787\,
            I => \N__34762\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__34786\,
            I => \N__34759\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__34785\,
            I => \N__34756\
        );

    \I__6256\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34751\
        );

    \I__6255\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34751\
        );

    \I__6254\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34744\
        );

    \I__6253\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34744\
        );

    \I__6252\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34744\
        );

    \I__6251\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34739\
        );

    \I__6250\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34739\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34736\
        );

    \I__6248\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34733\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34730\
        );

    \I__6246\ : InMux
    port map (
            O => \N__34762\,
            I => \N__34723\
        );

    \I__6245\ : InMux
    port map (
            O => \N__34759\,
            I => \N__34723\
        );

    \I__6244\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34723\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__34751\,
            I => \N__34718\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__34744\,
            I => \N__34718\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__34739\,
            I => eis_state_0
        );

    \I__6240\ : Odrv12
    port map (
            O => \N__34736\,
            I => eis_state_0
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__34733\,
            I => eis_state_0
        );

    \I__6238\ : Odrv12
    port map (
            O => \N__34730\,
            I => eis_state_0
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__34723\,
            I => eis_state_0
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__34718\,
            I => eis_state_0
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__34705\,
            I => \N__34702\
        );

    \I__6234\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34692\
        );

    \I__6233\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34687\
        );

    \I__6232\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34687\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__34699\,
            I => \N__34682\
        );

    \I__6230\ : CascadeMux
    port map (
            O => \N__34698\,
            I => \N__34679\
        );

    \I__6229\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34673\
        );

    \I__6228\ : InMux
    port map (
            O => \N__34696\,
            I => \N__34673\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__34695\,
            I => \N__34667\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34663\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34660\
        );

    \I__6224\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34655\
        );

    \I__6223\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34655\
        );

    \I__6222\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34648\
        );

    \I__6221\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34648\
        );

    \I__6220\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34648\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34645\
        );

    \I__6218\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34640\
        );

    \I__6217\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34640\
        );

    \I__6216\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34633\
        );

    \I__6215\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34633\
        );

    \I__6214\ : InMux
    port map (
            O => \N__34666\,
            I => \N__34633\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__34663\,
            I => eis_state_2
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__34660\,
            I => eis_state_2
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__34655\,
            I => eis_state_2
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__34648\,
            I => eis_state_2
        );

    \I__6209\ : Odrv4
    port map (
            O => \N__34645\,
            I => eis_state_2
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__34640\,
            I => eis_state_2
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__34633\,
            I => eis_state_2
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__34618\,
            I => \n12450_cascade_\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__34615\,
            I => \N__34611\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__34614\,
            I => \N__34608\
        );

    \I__6203\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34605\
        );

    \I__6202\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34602\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__34605\,
            I => \N__34599\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__34602\,
            I => \N__34596\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__34599\,
            I => \N__34593\
        );

    \I__6198\ : Span4Mux_h
    port map (
            O => \N__34596\,
            I => \N__34590\
        );

    \I__6197\ : Span4Mux_v
    port map (
            O => \N__34593\,
            I => \N__34586\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__34590\,
            I => \N__34583\
        );

    \I__6195\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34580\
        );

    \I__6194\ : Odrv4
    port map (
            O => \N__34586\,
            I => cmd_rdadctmp_16
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__34583\,
            I => cmd_rdadctmp_16
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__34580\,
            I => cmd_rdadctmp_16
        );

    \I__6191\ : SRMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__6189\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34564\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__34564\,
            I => n22120
        );

    \I__6187\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34558\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__34558\,
            I => n22312
        );

    \I__6185\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34552\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34552\,
            I => n23330
        );

    \I__6183\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34543\
        );

    \I__6182\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34543\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__34543\,
            I => n17633
        );

    \I__6180\ : SRMux
    port map (
            O => \N__34540\,
            I => \N__34537\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__34537\,
            I => \N__34531\
        );

    \I__6178\ : SRMux
    port map (
            O => \N__34536\,
            I => \N__34528\
        );

    \I__6177\ : SRMux
    port map (
            O => \N__34535\,
            I => \N__34525\
        );

    \I__6176\ : SRMux
    port map (
            O => \N__34534\,
            I => \N__34519\
        );

    \I__6175\ : Span4Mux_v
    port map (
            O => \N__34531\,
            I => \N__34511\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__34528\,
            I => \N__34511\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__34525\,
            I => \N__34511\
        );

    \I__6172\ : SRMux
    port map (
            O => \N__34524\,
            I => \N__34508\
        );

    \I__6171\ : SRMux
    port map (
            O => \N__34523\,
            I => \N__34505\
        );

    \I__6170\ : SRMux
    port map (
            O => \N__34522\,
            I => \N__34500\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34495\
        );

    \I__6168\ : SRMux
    port map (
            O => \N__34518\,
            I => \N__34492\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__34511\,
            I => \N__34485\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__34508\,
            I => \N__34485\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34485\
        );

    \I__6164\ : SRMux
    port map (
            O => \N__34504\,
            I => \N__34482\
        );

    \I__6163\ : SRMux
    port map (
            O => \N__34503\,
            I => \N__34479\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__34500\,
            I => \N__34476\
        );

    \I__6161\ : SRMux
    port map (
            O => \N__34499\,
            I => \N__34473\
        );

    \I__6160\ : SRMux
    port map (
            O => \N__34498\,
            I => \N__34470\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__34495\,
            I => \N__34465\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__34492\,
            I => \N__34465\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34458\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34458\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__34479\,
            I => \N__34458\
        );

    \I__6154\ : Span4Mux_v
    port map (
            O => \N__34476\,
            I => \N__34451\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34451\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__34470\,
            I => \N__34451\
        );

    \I__6151\ : Span4Mux_v
    port map (
            O => \N__34465\,
            I => \N__34448\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__34458\,
            I => \N__34443\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__34451\,
            I => \N__34443\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__34448\,
            I => \N__34440\
        );

    \I__6147\ : Span4Mux_h
    port map (
            O => \N__34443\,
            I => \N__34437\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__34440\,
            I => \N__34432\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__34437\,
            I => \N__34432\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__34432\,
            I => \iac_raw_buf_N_821\
        );

    \I__6143\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34426\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__34426\,
            I => n17_adj_1742
        );

    \I__6141\ : CEMux
    port map (
            O => \N__34423\,
            I => \N__34420\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34416\
        );

    \I__6139\ : CEMux
    port map (
            O => \N__34419\,
            I => \N__34413\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__34416\,
            I => \N__34410\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__34413\,
            I => \N__34405\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__34410\,
            I => \N__34405\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__34405\,
            I => n12369
        );

    \I__6134\ : CascadeMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__34393\,
            I => n24_adj_1503
        );

    \I__6130\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34382\
        );

    \I__6128\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34379\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__34385\,
            I => \N__34376\
        );

    \I__6126\ : Span12Mux_v
    port map (
            O => \N__34382\,
            I => \N__34373\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__34379\,
            I => \N__34370\
        );

    \I__6124\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34367\
        );

    \I__6123\ : Span12Mux_h
    port map (
            O => \N__34373\,
            I => \N__34364\
        );

    \I__6122\ : Span4Mux_h
    port map (
            O => \N__34370\,
            I => \N__34361\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__34367\,
            I => buf_adcdata_iac_16
        );

    \I__6120\ : Odrv12
    port map (
            O => \N__34364\,
            I => buf_adcdata_iac_16
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__34361\,
            I => buf_adcdata_iac_16
        );

    \I__6118\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34351\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__34351\,
            I => \N__34348\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__34348\,
            I => n23324
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__34345\,
            I => \N__34340\
        );

    \I__6114\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34335\
        );

    \I__6113\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34335\
        );

    \I__6112\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34332\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__34335\,
            I => req_data_cnt_8
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__34332\,
            I => req_data_cnt_8
        );

    \I__6109\ : CascadeMux
    port map (
            O => \N__34327\,
            I => \n19_adj_1727_cascade_\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__34324\,
            I => \n29_adj_1770_cascade_\
        );

    \I__6107\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34317\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__34320\,
            I => \N__34314\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34311\
        );

    \I__6104\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34308\
        );

    \I__6103\ : Span4Mux_v
    port map (
            O => \N__34311\,
            I => \N__34305\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__34308\,
            I => comm_test_buf_24_14
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__34305\,
            I => comm_test_buf_24_14
        );

    \I__6100\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34294\
        );

    \I__6099\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34294\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__34294\,
            I => \N__34290\
        );

    \I__6097\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34287\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__34290\,
            I => \N__34284\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34281\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__34284\,
            I => comm_test_buf_24_6
        );

    \I__6093\ : Odrv12
    port map (
            O => \N__34281\,
            I => comm_test_buf_24_6
        );

    \I__6092\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34271\
        );

    \I__6091\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34266\
        );

    \I__6090\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34266\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__34271\,
            I => n16_adj_1683
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__34266\,
            I => n16_adj_1683
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__34261\,
            I => \n17642_cascade_\
        );

    \I__6086\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34254\
        );

    \I__6085\ : InMux
    port map (
            O => \N__34257\,
            I => \N__34251\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__34254\,
            I => comm_test_buf_24_11
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34251\,
            I => comm_test_buf_24_11
        );

    \I__6082\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34240\
        );

    \I__6081\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34240\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__34240\,
            I => comm_test_buf_24_12
        );

    \I__6079\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34234\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__34231\,
            I => n13237
        );

    \I__6076\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34225\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__6074\ : Span4Mux_v
    port map (
            O => \N__34222\,
            I => \N__34219\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__34219\,
            I => n22295
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__34216\,
            I => \N__34213\
        );

    \I__6071\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34210\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__34207\,
            I => n4_adj_1667
        );

    \I__6068\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34201\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__34201\,
            I => \N__34198\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__34198\,
            I => n23294
        );

    \I__6065\ : InMux
    port map (
            O => \N__34195\,
            I => \N__34192\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__34192\,
            I => \N__34189\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__34189\,
            I => n30_adj_1588
        );

    \I__6062\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__34180\,
            I => \N__34175\
        );

    \I__6059\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34172\
        );

    \I__6058\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34169\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__34175\,
            I => comm_test_buf_24_3
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__34172\,
            I => comm_test_buf_24_3
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__34169\,
            I => comm_test_buf_24_3
        );

    \I__6054\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34159\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__34159\,
            I => n111_adj_1794
        );

    \I__6052\ : SRMux
    port map (
            O => \N__34156\,
            I => \N__34153\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34153\,
            I => n15545
        );

    \I__6050\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34147\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__34147\,
            I => \N__34144\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__34144\,
            I => \N__34140\
        );

    \I__6047\ : CascadeMux
    port map (
            O => \N__34143\,
            I => \N__34137\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__34140\,
            I => \N__34133\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34128\
        );

    \I__6044\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34128\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__34133\,
            I => buf_dds1_8
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__34128\,
            I => buf_dds1_8
        );

    \I__6041\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__34117\,
            I => n1_adj_1665
        );

    \I__6038\ : SRMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__6036\ : Span4Mux_h
    port map (
            O => \N__34108\,
            I => \N__34105\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__34105\,
            I => \comm_spi.data_tx_7__N_865\
        );

    \I__6034\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34095\
        );

    \I__6032\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34092\
        );

    \I__6031\ : Span4Mux_v
    port map (
            O => \N__34095\,
            I => \N__34088\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34085\
        );

    \I__6029\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34082\
        );

    \I__6028\ : Span4Mux_v
    port map (
            O => \N__34088\,
            I => \N__34077\
        );

    \I__6027\ : Span4Mux_h
    port map (
            O => \N__34085\,
            I => \N__34077\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__34082\,
            I => comm_test_buf_24_4
        );

    \I__6025\ : Odrv4
    port map (
            O => \N__34077\,
            I => comm_test_buf_24_4
        );

    \I__6024\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34069\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__34069\,
            I => n13231
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__34066\,
            I => \n19_adj_1710_cascade_\
        );

    \I__6021\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34060\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__34060\,
            I => \N__34057\
        );

    \I__6019\ : Span12Mux_h
    port map (
            O => \N__34057\,
            I => \N__34054\
        );

    \I__6018\ : Odrv12
    port map (
            O => \N__34054\,
            I => buf_data_iac_1
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__34051\,
            I => \n22_adj_1711_cascade_\
        );

    \I__6016\ : CascadeMux
    port map (
            O => \N__34048\,
            I => \n30_adj_1712_cascade_\
        );

    \I__6015\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34042\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__34042\,
            I => \N__34039\
        );

    \I__6013\ : Span4Mux_v
    port map (
            O => \N__34039\,
            I => \N__34036\
        );

    \I__6012\ : Span4Mux_v
    port map (
            O => \N__34036\,
            I => \N__34032\
        );

    \I__6011\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34029\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__34032\,
            I => \N__34024\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__34024\
        );

    \I__6008\ : Span4Mux_h
    port map (
            O => \N__34024\,
            I => \N__34020\
        );

    \I__6007\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34017\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__34020\,
            I => \comm_spi.n24031\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__34017\,
            I => \comm_spi.n24031\
        );

    \I__6004\ : InMux
    port map (
            O => \N__34012\,
            I => \N__34009\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__34009\,
            I => n30_adj_1705
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__34006\,
            I => \N__34003\
        );

    \I__6001\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33997\
        );

    \I__6000\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33994\
        );

    \I__5999\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33982\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__34000\,
            I => \N__33975\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__33997\,
            I => \N__33967\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__33994\,
            I => \N__33967\
        );

    \I__5995\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33962\
        );

    \I__5994\ : InMux
    port map (
            O => \N__33992\,
            I => \N__33962\
        );

    \I__5993\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33955\
        );

    \I__5992\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33955\
        );

    \I__5991\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33955\
        );

    \I__5990\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33945\
        );

    \I__5989\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33945\
        );

    \I__5988\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33940\
        );

    \I__5987\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33940\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__33982\,
            I => \N__33931\
        );

    \I__5985\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33928\
        );

    \I__5984\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33921\
        );

    \I__5983\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33921\
        );

    \I__5982\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33921\
        );

    \I__5981\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33914\
        );

    \I__5980\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33914\
        );

    \I__5979\ : InMux
    port map (
            O => \N__33973\,
            I => \N__33914\
        );

    \I__5978\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33911\
        );

    \I__5977\ : Span4Mux_v
    port map (
            O => \N__33967\,
            I => \N__33908\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__33962\,
            I => \N__33903\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__33955\,
            I => \N__33903\
        );

    \I__5974\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33897\
        );

    \I__5973\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33897\
        );

    \I__5972\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33892\
        );

    \I__5971\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33892\
        );

    \I__5970\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33889\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__33945\,
            I => \N__33886\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33883\
        );

    \I__5967\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33880\
        );

    \I__5966\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33877\
        );

    \I__5965\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33868\
        );

    \I__5964\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33868\
        );

    \I__5963\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33868\
        );

    \I__5962\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33868\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__33931\,
            I => \N__33861\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33861\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__33921\,
            I => \N__33861\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33858\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__33911\,
            I => \N__33851\
        );

    \I__5956\ : Span4Mux_h
    port map (
            O => \N__33908\,
            I => \N__33851\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__33903\,
            I => \N__33851\
        );

    \I__5954\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33848\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__33897\,
            I => \N__33845\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33836\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33836\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__33886\,
            I => \N__33836\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__33883\,
            I => \N__33836\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__33880\,
            I => \N__33823\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33823\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33823\
        );

    \I__5945\ : Span4Mux_v
    port map (
            O => \N__33861\,
            I => \N__33823\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__33858\,
            I => \N__33823\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__33851\,
            I => \N__33823\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33820\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__33845\,
            I => \N__33815\
        );

    \I__5940\ : Span4Mux_v
    port map (
            O => \N__33836\,
            I => \N__33815\
        );

    \I__5939\ : Span4Mux_h
    port map (
            O => \N__33823\,
            I => \N__33812\
        );

    \I__5938\ : Odrv12
    port map (
            O => \N__33820\,
            I => n13847
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__33815\,
            I => n13847
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__33812\,
            I => n13847
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__33805\,
            I => \N__33801\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__33804\,
            I => \N__33798\
        );

    \I__5933\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33794\
        );

    \I__5932\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33789\
        );

    \I__5931\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33789\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__33794\,
            I => cmd_rdadctmp_9_adj_1539
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__33789\,
            I => cmd_rdadctmp_9_adj_1539
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__33784\,
            I => \n2_adj_1666_cascade_\
        );

    \I__5927\ : SRMux
    port map (
            O => \N__33781\,
            I => \N__33778\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__33778\,
            I => \N__33775\
        );

    \I__5925\ : Odrv12
    port map (
            O => \N__33775\,
            I => \ADC_VDC.n17542\
        );

    \I__5924\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33768\
        );

    \I__5923\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33765\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__33768\,
            I => \N__33762\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33759\
        );

    \I__5920\ : Span4Mux_v
    port map (
            O => \N__33762\,
            I => \N__33756\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__33759\,
            I => \N__33753\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__33756\,
            I => \comm_spi.n15361\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__33753\,
            I => \comm_spi.n15361\
        );

    \I__5916\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33745\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__33745\,
            I => \N__33742\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__33742\,
            I => \N__33738\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__33741\,
            I => \N__33735\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__33738\,
            I => \N__33732\
        );

    \I__5911\ : InMux
    port map (
            O => \N__33735\,
            I => \N__33729\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__33732\,
            I => buf_adcdata_vdc_3
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__33729\,
            I => buf_adcdata_vdc_3
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__33724\,
            I => \n19_adj_1703_cascade_\
        );

    \I__5907\ : InMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__33718\,
            I => \N__33715\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__33715\,
            I => \N__33712\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__33712\,
            I => \N__33709\
        );

    \I__5903\ : Span4Mux_h
    port map (
            O => \N__33709\,
            I => \N__33706\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__33706\,
            I => buf_data_iac_3
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__33703\,
            I => \n22_adj_1704_cascade_\
        );

    \I__5900\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33697\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33694\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__33694\,
            I => \N__33691\
        );

    \I__5897\ : Sp12to4
    port map (
            O => \N__33691\,
            I => \N__33686\
        );

    \I__5896\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33681\
        );

    \I__5895\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33681\
        );

    \I__5894\ : Odrv12
    port map (
            O => \N__33686\,
            I => buf_adcdata_iac_3
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__33681\,
            I => buf_adcdata_iac_3
        );

    \I__5892\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33673\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__33673\,
            I => \N__33670\
        );

    \I__5890\ : Span12Mux_v
    port map (
            O => \N__33670\,
            I => \N__33665\
        );

    \I__5889\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33660\
        );

    \I__5888\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33660\
        );

    \I__5887\ : Odrv12
    port map (
            O => \N__33665\,
            I => cmd_rdadctmp_11_adj_1537
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__33660\,
            I => cmd_rdadctmp_11_adj_1537
        );

    \I__5885\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__5883\ : Span4Mux_v
    port map (
            O => \N__33649\,
            I => \N__33646\
        );

    \I__5882\ : Sp12to4
    port map (
            O => \N__33646\,
            I => \N__33641\
        );

    \I__5881\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33636\
        );

    \I__5880\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33636\
        );

    \I__5879\ : Odrv12
    port map (
            O => \N__33641\,
            I => buf_adcdata_vac_3
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__33636\,
            I => buf_adcdata_vac_3
        );

    \I__5877\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33628\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33624\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__33627\,
            I => \N__33621\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__33624\,
            I => \N__33618\
        );

    \I__5873\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33615\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__33618\,
            I => buf_adcdata_vdc_1
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__33615\,
            I => buf_adcdata_vdc_1
        );

    \I__5870\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33603\
        );

    \I__5868\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33599\
        );

    \I__5867\ : Span12Mux_h
    port map (
            O => \N__33603\,
            I => \N__33596\
        );

    \I__5866\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33593\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__33599\,
            I => buf_adcdata_vac_1
        );

    \I__5864\ : Odrv12
    port map (
            O => \N__33596\,
            I => buf_adcdata_vac_1
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__33593\,
            I => buf_adcdata_vac_1
        );

    \I__5862\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33570\
        );

    \I__5860\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33567\
        );

    \I__5859\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33564\
        );

    \I__5858\ : InMux
    port map (
            O => \N__33580\,
            I => \N__33561\
        );

    \I__5857\ : InMux
    port map (
            O => \N__33579\,
            I => \N__33556\
        );

    \I__5856\ : InMux
    port map (
            O => \N__33578\,
            I => \N__33556\
        );

    \I__5855\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33553\
        );

    \I__5854\ : InMux
    port map (
            O => \N__33576\,
            I => \N__33545\
        );

    \I__5853\ : InMux
    port map (
            O => \N__33575\,
            I => \N__33542\
        );

    \I__5852\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33537\
        );

    \I__5851\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33537\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__33570\,
            I => \N__33526\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__33567\,
            I => \N__33526\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__33564\,
            I => \N__33517\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__33561\,
            I => \N__33517\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__33556\,
            I => \N__33517\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__33553\,
            I => \N__33517\
        );

    \I__5844\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33513\
        );

    \I__5843\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33510\
        );

    \I__5842\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33507\
        );

    \I__5841\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33504\
        );

    \I__5840\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33501\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__33545\,
            I => \N__33494\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__33542\,
            I => \N__33494\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__33537\,
            I => \N__33494\
        );

    \I__5836\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33485\
        );

    \I__5835\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33485\
        );

    \I__5834\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33485\
        );

    \I__5833\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33485\
        );

    \I__5832\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33480\
        );

    \I__5831\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33480\
        );

    \I__5830\ : Span4Mux_v
    port map (
            O => \N__33526\,
            I => \N__33475\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__33517\,
            I => \N__33475\
        );

    \I__5828\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33472\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__33513\,
            I => \N__33467\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__33510\,
            I => \N__33467\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33507\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__33504\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__33501\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5822\ : Odrv12
    port map (
            O => \N__33494\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__33485\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__33480\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__33475\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__33472\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__33467\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__33448\,
            I => \N__33433\
        );

    \I__5815\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33426\
        );

    \I__5814\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33411\
        );

    \I__5813\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33411\
        );

    \I__5812\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33411\
        );

    \I__5811\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33411\
        );

    \I__5810\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33411\
        );

    \I__5809\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33411\
        );

    \I__5808\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33411\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__33439\,
            I => \N__33407\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__33438\,
            I => \N__33404\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__33437\,
            I => \N__33399\
        );

    \I__5804\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33388\
        );

    \I__5803\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33388\
        );

    \I__5802\ : CascadeMux
    port map (
            O => \N__33432\,
            I => \N__33382\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__33431\,
            I => \N__33375\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33372\
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__33429\,
            I => \N__33369\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33363\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__33411\,
            I => \N__33363\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33356\
        );

    \I__5795\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33356\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33356\
        );

    \I__5793\ : CascadeMux
    port map (
            O => \N__33403\,
            I => \N__33349\
        );

    \I__5792\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33333\
        );

    \I__5791\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33333\
        );

    \I__5790\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33333\
        );

    \I__5789\ : InMux
    port map (
            O => \N__33397\,
            I => \N__33333\
        );

    \I__5788\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33333\
        );

    \I__5787\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33333\
        );

    \I__5786\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33333\
        );

    \I__5785\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33330\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33327\
        );

    \I__5783\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33320\
        );

    \I__5782\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33320\
        );

    \I__5781\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33320\
        );

    \I__5780\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33315\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__33381\,
            I => \N__33311\
        );

    \I__5778\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33308\
        );

    \I__5777\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33303\
        );

    \I__5776\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33303\
        );

    \I__5775\ : InMux
    port map (
            O => \N__33375\,
            I => \N__33300\
        );

    \I__5774\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33295\
        );

    \I__5773\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33295\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__33368\,
            I => \N__33292\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__33363\,
            I => \N__33285\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33285\
        );

    \I__5769\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33274\
        );

    \I__5768\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33274\
        );

    \I__5767\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33274\
        );

    \I__5766\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33274\
        );

    \I__5765\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33274\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__33348\,
            I => \N__33270\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33267\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__33330\,
            I => \N__33261\
        );

    \I__5761\ : Span4Mux_h
    port map (
            O => \N__33327\,
            I => \N__33261\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__33320\,
            I => \N__33258\
        );

    \I__5759\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33253\
        );

    \I__5758\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33253\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__33315\,
            I => \N__33250\
        );

    \I__5756\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33246\
        );

    \I__5755\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33243\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33240\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33233\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__33300\,
            I => \N__33233\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__33295\,
            I => \N__33233\
        );

    \I__5750\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33226\
        );

    \I__5749\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33226\
        );

    \I__5748\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33226\
        );

    \I__5747\ : Span4Mux_v
    port map (
            O => \N__33285\,
            I => \N__33221\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33221\
        );

    \I__5745\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33218\
        );

    \I__5744\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33215\
        );

    \I__5743\ : Span12Mux_v
    port map (
            O => \N__33267\,
            I => \N__33212\
        );

    \I__5742\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33209\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__33261\,
            I => \N__33206\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__33258\,
            I => \N__33201\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33201\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__33250\,
            I => \N__33198\
        );

    \I__5737\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33195\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33182\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33182\
        );

    \I__5734\ : Span4Mux_h
    port map (
            O => \N__33240\,
            I => \N__33182\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__33233\,
            I => \N__33182\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__33226\,
            I => \N__33182\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__33221\,
            I => \N__33182\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__33218\,
            I => adc_state_2_adj_1550
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__33215\,
            I => adc_state_2_adj_1550
        );

    \I__5728\ : Odrv12
    port map (
            O => \N__33212\,
            I => adc_state_2_adj_1550
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__33209\,
            I => adc_state_2_adj_1550
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__33206\,
            I => adc_state_2_adj_1550
        );

    \I__5725\ : Odrv4
    port map (
            O => \N__33201\,
            I => adc_state_2_adj_1550
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__33198\,
            I => adc_state_2_adj_1550
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__33195\,
            I => adc_state_2_adj_1550
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__33182\,
            I => adc_state_2_adj_1550
        );

    \I__5721\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__33160\,
            I => \ADC_VDC.n11183\
        );

    \I__5719\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33154\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__33154\,
            I => \ADC_VDC.n23528\
        );

    \I__5717\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33147\
        );

    \I__5716\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33141\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__33147\,
            I => \N__33138\
        );

    \I__5714\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33135\
        );

    \I__5713\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33130\
        );

    \I__5712\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33130\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__33141\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__33138\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__33135\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__33130\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33121\,
            I => \bfn_11_6_0_\
        );

    \I__5706\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33112\
        );

    \I__5705\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33109\
        );

    \I__5704\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33106\
        );

    \I__5703\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33103\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33096\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__33109\,
            I => \N__33096\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33096\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__33103\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__33096\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33091\,
            I => \ADC_VDC.n20812\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__33088\,
            I => \N__33083\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__33087\,
            I => \N__33080\
        );

    \I__5694\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33077\
        );

    \I__5693\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33073\
        );

    \I__5692\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33070\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__33077\,
            I => \N__33067\
        );

    \I__5690\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33063\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33056\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33056\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__33067\,
            I => \N__33056\
        );

    \I__5686\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33053\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__33063\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__33056\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__33053\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__5682\ : InMux
    port map (
            O => \N__33046\,
            I => \ADC_VDC.n20813\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33036\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33033\
        );

    \I__5679\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33028\
        );

    \I__5678\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33028\
        );

    \I__5677\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33025\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33022\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__33033\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__33028\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__33025\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__33022\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__5671\ : InMux
    port map (
            O => \N__33013\,
            I => \ADC_VDC.n20814\
        );

    \I__5670\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33003\
        );

    \I__5669\ : InMux
    port map (
            O => \N__33009\,
            I => \N__33000\
        );

    \I__5668\ : InMux
    port map (
            O => \N__33008\,
            I => \N__32997\
        );

    \I__5667\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32992\
        );

    \I__5666\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32992\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__33003\,
            I => \N__32989\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__33000\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__32997\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__32992\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__32989\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__5660\ : InMux
    port map (
            O => \N__32980\,
            I => \ADC_VDC.n20815\
        );

    \I__5659\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32973\
        );

    \I__5658\ : InMux
    port map (
            O => \N__32976\,
            I => \N__32970\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__32973\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__32970\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__5655\ : InMux
    port map (
            O => \N__32965\,
            I => \ADC_VDC.n20816\
        );

    \I__5654\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32958\
        );

    \I__5653\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32955\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__32958\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__32955\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__5650\ : InMux
    port map (
            O => \N__32950\,
            I => \ADC_VDC.n20817\
        );

    \I__5649\ : InMux
    port map (
            O => \N__32947\,
            I => \ADC_VDC.n20818\
        );

    \I__5648\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32940\
        );

    \I__5647\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32937\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__32940\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__32937\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__5644\ : CEMux
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32926\
        );

    \I__5642\ : Odrv12
    port map (
            O => \N__32926\,
            I => \ADC_VDC.n17565\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__5640\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32914\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__32914\,
            I => \SIG_DDS.tmp_buf_10\
        );

    \I__5637\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__32908\,
            I => \N__32905\
        );

    \I__5635\ : Span12Mux_v
    port map (
            O => \N__32905\,
            I => \N__32900\
        );

    \I__5634\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32897\
        );

    \I__5633\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32894\
        );

    \I__5632\ : Odrv12
    port map (
            O => \N__32900\,
            I => buf_dds0_11
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__32897\,
            I => buf_dds0_11
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__32894\,
            I => buf_dds0_11
        );

    \I__5629\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32884\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__32884\,
            I => \SIG_DDS.tmp_buf_11\
        );

    \I__5627\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32878\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__32878\,
            I => \ADC_VDC.n22063\
        );

    \I__5625\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32869\
        );

    \I__5624\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32862\
        );

    \I__5623\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32862\
        );

    \I__5622\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32862\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__32869\,
            I => \N__32857\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32857\
        );

    \I__5619\ : Odrv12
    port map (
            O => \N__32857\,
            I => \RTD.n20050\
        );

    \I__5618\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32845\
        );

    \I__5617\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32840\
        );

    \I__5616\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32840\
        );

    \I__5615\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32837\
        );

    \I__5614\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32834\
        );

    \I__5613\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32830\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__32848\,
            I => \N__32825\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__32845\,
            I => \N__32820\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32820\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32815\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__32834\,
            I => \N__32815\
        );

    \I__5607\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32812\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__32830\,
            I => \N__32809\
        );

    \I__5605\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32804\
        );

    \I__5604\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32804\
        );

    \I__5603\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32801\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__32820\,
            I => \N__32795\
        );

    \I__5601\ : Span4Mux_v
    port map (
            O => \N__32815\,
            I => \N__32795\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32792\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__32809\,
            I => \N__32785\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32785\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32785\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__32800\,
            I => \N__32782\
        );

    \I__5595\ : Span4Mux_v
    port map (
            O => \N__32795\,
            I => \N__32779\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__32792\,
            I => \N__32774\
        );

    \I__5593\ : Span4Mux_v
    port map (
            O => \N__32785\,
            I => \N__32774\
        );

    \I__5592\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32771\
        );

    \I__5591\ : Sp12to4
    port map (
            O => \N__32779\,
            I => \N__32768\
        );

    \I__5590\ : Span4Mux_v
    port map (
            O => \N__32774\,
            I => \N__32765\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__32771\,
            I => \N__32762\
        );

    \I__5588\ : Span12Mux_h
    port map (
            O => \N__32768\,
            I => \N__32755\
        );

    \I__5587\ : Sp12to4
    port map (
            O => \N__32765\,
            I => \N__32755\
        );

    \I__5586\ : Span12Mux_v
    port map (
            O => \N__32762\,
            I => \N__32755\
        );

    \I__5585\ : Odrv12
    port map (
            O => \N__32755\,
            I => \VDC_SDO\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__32752\,
            I => \ADC_VDC.n35_cascade_\
        );

    \I__5583\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32746\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__32746\,
            I => \ADC_VDC.n45\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__32743\,
            I => \N__32740\
        );

    \I__5580\ : InMux
    port map (
            O => \N__32740\,
            I => \N__32737\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__32737\,
            I => \ADC_VDC.n22067\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__32734\,
            I => \N__32719\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__32733\,
            I => \N__32716\
        );

    \I__5576\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32704\
        );

    \I__5575\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32697\
        );

    \I__5574\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32689\
        );

    \I__5573\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32689\
        );

    \I__5572\ : InMux
    port map (
            O => \N__32728\,
            I => \N__32689\
        );

    \I__5571\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32679\
        );

    \I__5570\ : InMux
    port map (
            O => \N__32726\,
            I => \N__32679\
        );

    \I__5569\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32679\
        );

    \I__5568\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32679\
        );

    \I__5567\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32674\
        );

    \I__5566\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32674\
        );

    \I__5565\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32665\
        );

    \I__5564\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32665\
        );

    \I__5563\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32665\
        );

    \I__5562\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32665\
        );

    \I__5561\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32650\
        );

    \I__5560\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32650\
        );

    \I__5559\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32650\
        );

    \I__5558\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32650\
        );

    \I__5557\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32650\
        );

    \I__5556\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32650\
        );

    \I__5555\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32650\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__32704\,
            I => \N__32647\
        );

    \I__5553\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32642\
        );

    \I__5552\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32642\
        );

    \I__5551\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32638\
        );

    \I__5550\ : InMux
    port map (
            O => \N__32700\,
            I => \N__32635\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__32697\,
            I => \N__32632\
        );

    \I__5548\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32629\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32626\
        );

    \I__5546\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32623\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__32679\,
            I => \N__32608\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__32674\,
            I => \N__32608\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__32665\,
            I => \N__32608\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__32650\,
            I => \N__32608\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__32647\,
            I => \N__32600\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__32642\,
            I => \N__32600\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__32641\,
            I => \N__32592\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32577\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32577\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__32632\,
            I => \N__32577\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__32629\,
            I => \N__32577\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__32626\,
            I => \N__32577\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32577\
        );

    \I__5532\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32564\
        );

    \I__5531\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32564\
        );

    \I__5530\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32564\
        );

    \I__5529\ : InMux
    port map (
            O => \N__32619\,
            I => \N__32564\
        );

    \I__5528\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32564\
        );

    \I__5527\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32564\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__32608\,
            I => \N__32561\
        );

    \I__5525\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32556\
        );

    \I__5524\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32556\
        );

    \I__5523\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32553\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__32600\,
            I => \N__32550\
        );

    \I__5521\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32543\
        );

    \I__5520\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32543\
        );

    \I__5519\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32543\
        );

    \I__5518\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32536\
        );

    \I__5517\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32536\
        );

    \I__5516\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32536\
        );

    \I__5515\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32531\
        );

    \I__5514\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32531\
        );

    \I__5513\ : Span4Mux_v
    port map (
            O => \N__32577\,
            I => \N__32528\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__32564\,
            I => adc_state_3
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__32561\,
            I => adc_state_3
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__32556\,
            I => adc_state_3
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__32553\,
            I => adc_state_3
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__32550\,
            I => adc_state_3
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__32543\,
            I => adc_state_3
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__32536\,
            I => adc_state_3
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__32531\,
            I => adc_state_3
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__32528\,
            I => adc_state_3
        );

    \I__5503\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32498\
        );

    \I__5502\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32498\
        );

    \I__5501\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32498\
        );

    \I__5500\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32491\
        );

    \I__5499\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32487\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__32498\,
            I => \N__32481\
        );

    \I__5497\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32478\
        );

    \I__5496\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32473\
        );

    \I__5495\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32473\
        );

    \I__5494\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32467\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32464\
        );

    \I__5492\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32461\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__32487\,
            I => \N__32454\
        );

    \I__5490\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32451\
        );

    \I__5489\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32447\
        );

    \I__5488\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32444\
        );

    \I__5487\ : Sp12to4
    port map (
            O => \N__32481\,
            I => \N__32441\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32438\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32435\
        );

    \I__5484\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32428\
        );

    \I__5483\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32428\
        );

    \I__5482\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32428\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__32467\,
            I => \N__32421\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__32464\,
            I => \N__32421\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32421\
        );

    \I__5478\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32414\
        );

    \I__5477\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32414\
        );

    \I__5476\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32414\
        );

    \I__5475\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32411\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__32454\,
            I => \N__32406\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32406\
        );

    \I__5472\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32403\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__32447\,
            I => adc_state_1_adj_1551
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32444\,
            I => adc_state_1_adj_1551
        );

    \I__5469\ : Odrv12
    port map (
            O => \N__32441\,
            I => adc_state_1_adj_1551
        );

    \I__5468\ : Odrv4
    port map (
            O => \N__32438\,
            I => adc_state_1_adj_1551
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__32435\,
            I => adc_state_1_adj_1551
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__32428\,
            I => adc_state_1_adj_1551
        );

    \I__5465\ : Odrv4
    port map (
            O => \N__32421\,
            I => adc_state_1_adj_1551
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__32414\,
            I => adc_state_1_adj_1551
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32411\,
            I => adc_state_1_adj_1551
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__32406\,
            I => adc_state_1_adj_1551
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__32403\,
            I => adc_state_1_adj_1551
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__32380\,
            I => \N__32377\
        );

    \I__5459\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32373\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__32376\,
            I => \N__32369\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32366\
        );

    \I__5456\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32363\
        );

    \I__5455\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32360\
        );

    \I__5454\ : Span4Mux_v
    port map (
            O => \N__32366\,
            I => \N__32357\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32354\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__32360\,
            I => buf_dds0_5
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__32357\,
            I => buf_dds0_5
        );

    \I__5450\ : Odrv12
    port map (
            O => \N__32354\,
            I => buf_dds0_5
        );

    \I__5449\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32344\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__32344\,
            I => \SIG_DDS.tmp_buf_4\
        );

    \I__5447\ : CascadeMux
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__5446\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32335\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__32335\,
            I => \SIG_DDS.tmp_buf_5\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__32332\,
            I => \N__32329\
        );

    \I__5443\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32326\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__32326\,
            I => \SIG_DDS.tmp_buf_9\
        );

    \I__5441\ : CascadeMux
    port map (
            O => \N__32323\,
            I => \N__32320\
        );

    \I__5440\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32317\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__32317\,
            I => \SIG_DDS.tmp_buf_6\
        );

    \I__5438\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32309\
        );

    \I__5437\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32306\
        );

    \I__5436\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32303\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32300\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__32306\,
            I => buf_dds0_7
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__32303\,
            I => buf_dds0_7
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__32300\,
            I => buf_dds0_7
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__32293\,
            I => \N__32290\
        );

    \I__5430\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32287\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32284\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__32284\,
            I => \N__32279\
        );

    \I__5427\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32276\
        );

    \I__5426\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32273\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__32279\,
            I => \N__32270\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32267\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__32273\,
            I => buf_dds0_12
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__32270\,
            I => buf_dds0_12
        );

    \I__5421\ : Odrv4
    port map (
            O => \N__32267\,
            I => buf_dds0_12
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__32260\,
            I => \N__32257\
        );

    \I__5419\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32254\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__32254\,
            I => \SIG_DDS.tmp_buf_12\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__32251\,
            I => \N__32248\
        );

    \I__5416\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32245\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__32245\,
            I => \SIG_DDS.tmp_buf_13\
        );

    \I__5414\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32239\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32236\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__32236\,
            I => \N__32232\
        );

    \I__5411\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32228\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__32232\,
            I => \N__32225\
        );

    \I__5409\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32222\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32219\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__32225\,
            I => buf_dds0_14
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__32222\,
            I => buf_dds0_14
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__32219\,
            I => buf_dds0_14
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__32212\,
            I => \N__32209\
        );

    \I__5403\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32206\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__32206\,
            I => \SIG_DDS.tmp_buf_14\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__32203\,
            I => \N__32200\
        );

    \I__5400\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32197\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__32197\,
            I => \N__32192\
        );

    \I__5398\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32189\
        );

    \I__5397\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32186\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__32192\,
            I => \N__32183\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__32189\,
            I => buf_dds0_15
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__32186\,
            I => buf_dds0_15
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__32183\,
            I => buf_dds0_15
        );

    \I__5392\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32173\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__32173\,
            I => \SIG_DDS.tmp_buf_7\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \N__32167\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32164\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__32164\,
            I => \SIG_DDS.tmp_buf_8\
        );

    \I__5387\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32157\
        );

    \I__5386\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32154\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__32157\,
            I => cmd_rdadctmp_6
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__32154\,
            I => cmd_rdadctmp_6
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__32149\,
            I => \N__32143\
        );

    \I__5382\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32137\
        );

    \I__5381\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32137\
        );

    \I__5380\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32132\
        );

    \I__5379\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32132\
        );

    \I__5378\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32129\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__32137\,
            I => acadc_dtrig_i
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32132\,
            I => acadc_dtrig_i
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__32129\,
            I => acadc_dtrig_i
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__32122\,
            I => \N__32118\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__32121\,
            I => \N__32115\
        );

    \I__5372\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32109\
        );

    \I__5371\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32109\
        );

    \I__5370\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32106\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__32109\,
            I => cmd_rdadctmp_29
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__32106\,
            I => cmd_rdadctmp_29
        );

    \I__5367\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32096\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__32100\,
            I => \N__32086\
        );

    \I__5365\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32083\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32080\
        );

    \I__5363\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32073\
        );

    \I__5362\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32073\
        );

    \I__5361\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32073\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__32092\,
            I => \N__32068\
        );

    \I__5359\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32061\
        );

    \I__5358\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32061\
        );

    \I__5357\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32056\
        );

    \I__5356\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32056\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__32083\,
            I => \N__32053\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__32080\,
            I => \N__32050\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32047\
        );

    \I__5352\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32044\
        );

    \I__5351\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32039\
        );

    \I__5350\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32039\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32034\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32034\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32029\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__32029\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__32053\,
            I => \N__32020\
        );

    \I__5344\ : Span4Mux_h
    port map (
            O => \N__32050\,
            I => \N__32020\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__32047\,
            I => \N__32020\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__32020\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__32039\,
            I => \DTRIG_N_1182_adj_1549\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__32034\,
            I => \DTRIG_N_1182_adj_1549\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__32029\,
            I => \DTRIG_N_1182_adj_1549\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__32020\,
            I => \DTRIG_N_1182_adj_1549\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__32011\,
            I => \N__32008\
        );

    \I__5336\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32005\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__32005\,
            I => \N__32001\
        );

    \I__5334\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31993\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__32001\,
            I => \N__31988\
        );

    \I__5332\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31981\
        );

    \I__5331\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31981\
        );

    \I__5330\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31981\
        );

    \I__5329\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31976\
        );

    \I__5328\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31976\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__31993\,
            I => \N__31973\
        );

    \I__5326\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31967\
        );

    \I__5325\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31964\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__31988\,
            I => \N__31958\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31958\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31953\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__31973\,
            I => \N__31953\
        );

    \I__5320\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31948\
        );

    \I__5319\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31948\
        );

    \I__5318\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31945\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31940\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__31964\,
            I => \N__31940\
        );

    \I__5315\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31937\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__31958\,
            I => \N__31934\
        );

    \I__5313\ : Span4Mux_h
    port map (
            O => \N__31953\,
            I => \N__31931\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__31948\,
            I => adc_state_1_adj_1515
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__31945\,
            I => adc_state_1_adj_1515
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__31940\,
            I => adc_state_1_adj_1515
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__31937\,
            I => adc_state_1_adj_1515
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__31934\,
            I => adc_state_1_adj_1515
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__31931\,
            I => adc_state_1_adj_1515
        );

    \I__5306\ : CascadeMux
    port map (
            O => \N__31918\,
            I => \N__31915\
        );

    \I__5305\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31906\
        );

    \I__5304\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31906\
        );

    \I__5303\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31901\
        );

    \I__5302\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31901\
        );

    \I__5301\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31898\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__31906\,
            I => acadc_dtrig_v
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__31901\,
            I => acadc_dtrig_v
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__31898\,
            I => acadc_dtrig_v
        );

    \I__5297\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31887\
        );

    \I__5296\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31884\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31881\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__31884\,
            I => \N__31878\
        );

    \I__5293\ : Span4Mux_h
    port map (
            O => \N__31881\,
            I => \N__31872\
        );

    \I__5292\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31872\
        );

    \I__5291\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31869\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__31872\,
            I => \N__31866\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__31869\,
            I => buf_dds1_9
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__31866\,
            I => buf_dds1_9
        );

    \I__5287\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31858\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__31858\,
            I => n23534
        );

    \I__5285\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31850\
        );

    \I__5284\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31845\
        );

    \I__5283\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31845\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__31850\,
            I => buf_dds0_10
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__31845\,
            I => buf_dds0_10
        );

    \I__5280\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31836\
        );

    \I__5279\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31833\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31830\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__31833\,
            I => \N__31826\
        );

    \I__5276\ : Span4Mux_v
    port map (
            O => \N__31830\,
            I => \N__31823\
        );

    \I__5275\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31820\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__31826\,
            I => \N__31817\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__31823\,
            I => buf_dds0_6
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__31820\,
            I => buf_dds0_6
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__31817\,
            I => buf_dds0_6
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__31810\,
            I => \n13_cascade_\
        );

    \I__5269\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31804\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__31804\,
            I => n22395
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__31801\,
            I => \N__31798\
        );

    \I__5266\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31794\
        );

    \I__5265\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31791\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31788\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31785\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__31788\,
            I => \N__31782\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__31785\,
            I => \N__31779\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__31782\,
            I => \N__31775\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__31779\,
            I => \N__31772\
        );

    \I__5258\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31769\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__31775\,
            I => cmd_rdadctmp_30
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__31772\,
            I => cmd_rdadctmp_30
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__31769\,
            I => cmd_rdadctmp_30
        );

    \I__5254\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31758\
        );

    \I__5253\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31755\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31752\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__31755\,
            I => n13_adj_1591
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__31752\,
            I => n13_adj_1591
        );

    \I__5249\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31744\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__31744\,
            I => n11_adj_1592
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__31741\,
            I => \n23510_cascade_\
        );

    \I__5246\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31732\
        );

    \I__5244\ : Odrv12
    port map (
            O => \N__31732\,
            I => n22276
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__31729\,
            I => \n23513_cascade_\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__31726\,
            I => \n30_adj_1759_cascade_\
        );

    \I__5241\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31720\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__31720\,
            I => n26_adj_1758
        );

    \I__5239\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31711\
        );

    \I__5238\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31711\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__31711\,
            I => eis_end
        );

    \I__5236\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31705\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__31705\,
            I => n112_adj_1762
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__31702\,
            I => \n21946_cascade_\
        );

    \I__5233\ : InMux
    port map (
            O => \N__31699\,
            I => \N__31696\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__31696\,
            I => n21880
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__31693\,
            I => \n24_cascade_\
        );

    \I__5230\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31687\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__31687\,
            I => \N__31684\
        );

    \I__5228\ : Span12Mux_s8_v
    port map (
            O => \N__31684\,
            I => \N__31680\
        );

    \I__5227\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31677\
        );

    \I__5226\ : Span12Mux_h
    port map (
            O => \N__31680\,
            I => \N__31673\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31670\
        );

    \I__5224\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31667\
        );

    \I__5223\ : Span12Mux_v
    port map (
            O => \N__31673\,
            I => \N__31664\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__31670\,
            I => \N__31661\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__31667\,
            I => buf_adcdata_iac_22
        );

    \I__5220\ : Odrv12
    port map (
            O => \N__31664\,
            I => buf_adcdata_iac_22
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__31661\,
            I => buf_adcdata_iac_22
        );

    \I__5218\ : IoInMux
    port map (
            O => \N__31654\,
            I => \N__31651\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31648\
        );

    \I__5216\ : Span12Mux_s1_h
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__5215\ : Span12Mux_h
    port map (
            O => \N__31645\,
            I => \N__31640\
        );

    \I__5214\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31635\
        );

    \I__5213\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31635\
        );

    \I__5212\ : Odrv12
    port map (
            O => \N__31640\,
            I => \VAC_FLT0\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__31635\,
            I => \VAC_FLT0\
        );

    \I__5210\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31627\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__31627\,
            I => \N__31624\
        );

    \I__5208\ : Odrv4
    port map (
            O => \N__31624\,
            I => n17_adj_1764
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__31621\,
            I => \n11981_cascade_\
        );

    \I__5206\ : IoInMux
    port map (
            O => \N__31618\,
            I => \N__31615\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__5204\ : IoSpan4Mux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__5203\ : Span4Mux_s3_h
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__31603\,
            I => \N__31599\
        );

    \I__5200\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31596\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__31599\,
            I => \N__31590\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__31596\,
            I => \N__31590\
        );

    \I__5197\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31587\
        );

    \I__5196\ : Span4Mux_v
    port map (
            O => \N__31590\,
            I => \N__31584\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__31587\,
            I => \VAC_FLT1\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__31584\,
            I => \VAC_FLT1\
        );

    \I__5193\ : InMux
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__31576\,
            I => n24_adj_1576
        );

    \I__5191\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31570\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__31570\,
            I => n11986
        );

    \I__5189\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31564\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31561\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__31561\,
            I => \N__31558\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__31558\,
            I => n30_adj_1692
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__31555\,
            I => \N__31552\
        );

    \I__5184\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31548\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__31551\,
            I => \N__31544\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__31548\,
            I => \N__31541\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__31547\,
            I => \N__31538\
        );

    \I__5180\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31535\
        );

    \I__5179\ : Span4Mux_h
    port map (
            O => \N__31541\,
            I => \N__31532\
        );

    \I__5178\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31529\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31526\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__31532\,
            I => \N__31523\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__31529\,
            I => cmd_rdadctmp_25_adj_1523
        );

    \I__5174\ : Odrv12
    port map (
            O => \N__31526\,
            I => cmd_rdadctmp_25_adj_1523
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__31523\,
            I => cmd_rdadctmp_25_adj_1523
        );

    \I__5172\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31513\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31509\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__31512\,
            I => \N__31506\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__31509\,
            I => \N__31503\
        );

    \I__5168\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31500\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__31503\,
            I => buf_adcdata_vdc_18
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__31500\,
            I => buf_adcdata_vdc_18
        );

    \I__5165\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__31492\,
            I => \N__31489\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5162\ : Sp12to4
    port map (
            O => \N__31486\,
            I => \N__31481\
        );

    \I__5161\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31478\
        );

    \I__5160\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31475\
        );

    \I__5159\ : Span12Mux_h
    port map (
            O => \N__31481\,
            I => \N__31472\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__31478\,
            I => \N__31469\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__31475\,
            I => buf_adcdata_vac_18
        );

    \I__5156\ : Odrv12
    port map (
            O => \N__31472\,
            I => buf_adcdata_vac_18
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__31469\,
            I => buf_adcdata_vac_18
        );

    \I__5154\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__31459\,
            I => n22163
        );

    \I__5152\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__31453\,
            I => \N__31449\
        );

    \I__5150\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31446\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__31449\,
            I => \comm_spi.n15360\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__31446\,
            I => \comm_spi.n15360\
        );

    \I__5147\ : SRMux
    port map (
            O => \N__31441\,
            I => \N__31438\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__31438\,
            I => \N__31435\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__31435\,
            I => \comm_spi.data_tx_7__N_857\
        );

    \I__5144\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31428\
        );

    \I__5143\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31425\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__31425\,
            I => comm_test_buf_24_19
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__31422\,
            I => comm_test_buf_24_19
        );

    \I__5139\ : InMux
    port map (
            O => \N__31417\,
            I => \N__31413\
        );

    \I__5138\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31410\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__31413\,
            I => comm_test_buf_24_20
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__31410\,
            I => comm_test_buf_24_20
        );

    \I__5135\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31402\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__31402\,
            I => \N__31399\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__31399\,
            I => \N__31396\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__31396\,
            I => n111_adj_1785
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__31393\,
            I => \N__31390\
        );

    \I__5130\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31384\
        );

    \I__5129\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31384\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__31384\,
            I => cmd_rdadctmp_7_adj_1541
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__31381\,
            I => \N__31378\
        );

    \I__5126\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31372\
        );

    \I__5125\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31372\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__31372\,
            I => cmd_rdadctmp_6_adj_1542
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__31369\,
            I => \N__31366\
        );

    \I__5122\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31360\
        );

    \I__5121\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31360\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__31360\,
            I => cmd_rdadctmp_5_adj_1543
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__31357\,
            I => \N__31353\
        );

    \I__5118\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31350\
        );

    \I__5117\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31347\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__31350\,
            I => \N__31344\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__31347\,
            I => cmd_rdadctmp_3_adj_1545
        );

    \I__5114\ : Odrv12
    port map (
            O => \N__31344\,
            I => cmd_rdadctmp_3_adj_1545
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__31339\,
            I => \N__31336\
        );

    \I__5112\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31330\
        );

    \I__5111\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31330\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__31330\,
            I => cmd_rdadctmp_4_adj_1544
        );

    \I__5109\ : InMux
    port map (
            O => \N__31327\,
            I => \N__31324\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__31324\,
            I => \N__31319\
        );

    \I__5107\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31316\
        );

    \I__5106\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31313\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__31319\,
            I => \N__31310\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__31316\,
            I => \N__31307\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__31313\,
            I => buf_dds1_6
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__31310\,
            I => buf_dds1_6
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__31307\,
            I => buf_dds1_6
        );

    \I__5100\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31297\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31294\
        );

    \I__5098\ : Span4Mux_v
    port map (
            O => \N__31294\,
            I => \N__31291\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__31291\,
            I => \N__31288\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__31288\,
            I => \N__31285\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__31285\,
            I => buf_data_iac_0
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__31282\,
            I => \N__31279\
        );

    \I__5093\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31276\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31272\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__31275\,
            I => \N__31269\
        );

    \I__5090\ : Span12Mux_v
    port map (
            O => \N__31272\,
            I => \N__31265\
        );

    \I__5089\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31262\
        );

    \I__5088\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31259\
        );

    \I__5087\ : Odrv12
    port map (
            O => \N__31265\,
            I => cmd_rdadctmp_21_adj_1527
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__31262\,
            I => cmd_rdadctmp_21_adj_1527
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__31259\,
            I => cmd_rdadctmp_21_adj_1527
        );

    \I__5084\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31248\
        );

    \I__5083\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31245\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__31248\,
            I => \N__31240\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31240\
        );

    \I__5080\ : Span4Mux_h
    port map (
            O => \N__31240\,
            I => \N__31237\
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__31237\,
            I => \comm_spi.n15369\
        );

    \I__5078\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31231\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__31231\,
            I => \N__31228\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__31228\,
            I => \N__31224\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__31227\,
            I => \N__31221\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__31224\,
            I => \N__31218\
        );

    \I__5073\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31215\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__31218\,
            I => \buf_readRTD_13\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__31215\,
            I => \buf_readRTD_13\
        );

    \I__5070\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31207\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__31204\,
            I => \N__31201\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__31201\,
            I => \N__31198\
        );

    \I__5066\ : Sp12to4
    port map (
            O => \N__31198\,
            I => \N__31193\
        );

    \I__5065\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31190\
        );

    \I__5064\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31187\
        );

    \I__5063\ : Span12Mux_h
    port map (
            O => \N__31193\,
            I => \N__31182\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__31190\,
            I => \N__31182\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__31187\,
            I => buf_adcdata_vac_21
        );

    \I__5060\ : Odrv12
    port map (
            O => \N__31182\,
            I => buf_adcdata_vac_21
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31174\
        );

    \I__5058\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31171\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__31171\,
            I => \N__31166\
        );

    \I__5056\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31163\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__31169\,
            I => \N__31160\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__31166\,
            I => \N__31153\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31153\
        );

    \I__5052\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31148\
        );

    \I__5051\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31148\
        );

    \I__5050\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31145\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__31153\,
            I => \N__31142\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__31148\,
            I => \buf_cfgRTD_5\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__31145\,
            I => \buf_cfgRTD_5\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__31142\,
            I => \buf_cfgRTD_5\
        );

    \I__5045\ : CascadeMux
    port map (
            O => \N__31135\,
            I => \n23384_cascade_\
        );

    \I__5044\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31129\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__31129\,
            I => \N__31126\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__31126\,
            I => \N__31122\
        );

    \I__5041\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31119\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__31122\,
            I => cmd_rdadcbuf_32
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__31119\,
            I => cmd_rdadcbuf_32
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__31114\,
            I => \N__31110\
        );

    \I__5037\ : CascadeMux
    port map (
            O => \N__31113\,
            I => \N__31107\
        );

    \I__5036\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31102\
        );

    \I__5035\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31102\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__31102\,
            I => buf_adcdata_vdc_21
        );

    \I__5033\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31096\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__31096\,
            I => \N__31092\
        );

    \I__5031\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__5030\ : Odrv12
    port map (
            O => \N__31092\,
            I => cmd_rdadcbuf_24
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__31089\,
            I => cmd_rdadcbuf_24
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__31084\,
            I => \N__31069\
        );

    \I__5027\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31057\
        );

    \I__5026\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31054\
        );

    \I__5025\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31037\
        );

    \I__5024\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31037\
        );

    \I__5023\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31037\
        );

    \I__5022\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31037\
        );

    \I__5021\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31037\
        );

    \I__5020\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31037\
        );

    \I__5019\ : InMux
    port map (
            O => \N__31075\,
            I => \N__31037\
        );

    \I__5018\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31037\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__31073\,
            I => \N__31034\
        );

    \I__5016\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31017\
        );

    \I__5015\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31017\
        );

    \I__5014\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31017\
        );

    \I__5013\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31017\
        );

    \I__5012\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31017\
        );

    \I__5011\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31017\
        );

    \I__5010\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31017\
        );

    \I__5009\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31008\
        );

    \I__5008\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31008\
        );

    \I__5007\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31008\
        );

    \I__5006\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31008\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__31057\,
            I => \N__31005\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31002\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__31037\,
            I => \N__30999\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31034\,
            I => \N__30996\
        );

    \I__5001\ : InMux
    port map (
            O => \N__31033\,
            I => \N__30991\
        );

    \I__5000\ : InMux
    port map (
            O => \N__31032\,
            I => \N__30991\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__30988\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__30985\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__31005\,
            I => \N__30982\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__31002\,
            I => \N__30977\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30977\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__30996\,
            I => n12352
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__30991\,
            I => n12352
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__30988\,
            I => n12352
        );

    \I__4991\ : Odrv12
    port map (
            O => \N__30985\,
            I => n12352
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__30982\,
            I => n12352
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__30977\,
            I => n12352
        );

    \I__4988\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30961\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30958\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__30958\,
            I => \N__30954\
        );

    \I__4985\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30951\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__30954\,
            I => cmd_rdadcbuf_11
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__30951\,
            I => cmd_rdadcbuf_11
        );

    \I__4982\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30942\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__30945\,
            I => \N__30939\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30936\
        );

    \I__4979\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30933\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__30936\,
            I => buf_adcdata_vdc_12
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__30933\,
            I => buf_adcdata_vdc_12
        );

    \I__4976\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30925\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30922\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__30922\,
            I => \N__30919\
        );

    \I__4973\ : Span4Mux_h
    port map (
            O => \N__30919\,
            I => \N__30915\
        );

    \I__4972\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30912\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__30915\,
            I => \N__30908\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30905\
        );

    \I__4969\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30902\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__30908\,
            I => \N__30899\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__30905\,
            I => \N__30896\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__30902\,
            I => buf_adcdata_vac_12
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__30899\,
            I => buf_adcdata_vac_12
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__30896\,
            I => buf_adcdata_vac_12
        );

    \I__4963\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30886\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30883\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__30883\,
            I => \N__30879\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__30882\,
            I => \N__30876\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__30879\,
            I => \N__30873\
        );

    \I__4958\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30870\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__30873\,
            I => \buf_readRTD_4\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__30870\,
            I => \buf_readRTD_4\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__30865\,
            I => \n19_adj_1734_cascade_\
        );

    \I__4954\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30859\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__4952\ : Span4Mux_v
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__30853\,
            I => \ADC_VDC.n21991\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \ADC_VDC.n22075_cascade_\
        );

    \I__4949\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30844\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__30844\,
            I => \ADC_VDC.n44_adj_1487\
        );

    \I__4947\ : CEMux
    port map (
            O => \N__30841\,
            I => \N__30838\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30835\
        );

    \I__4945\ : Odrv12
    port map (
            O => \N__30835\,
            I => \ADC_VDC.n39_adj_1488\
        );

    \I__4944\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30829\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__30829\,
            I => \ADC_VDC.n6_adj_1485\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__30826\,
            I => \ADC_VDC.n21859_cascade_\
        );

    \I__4941\ : CascadeMux
    port map (
            O => \N__30823\,
            I => \ADC_VDC.n22628_cascade_\
        );

    \I__4940\ : InMux
    port map (
            O => \N__30820\,
            I => \N__30816\
        );

    \I__4939\ : InMux
    port map (
            O => \N__30819\,
            I => \N__30813\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__30816\,
            I => \ADC_VDC.n21859\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__30813\,
            I => \ADC_VDC.n21859\
        );

    \I__4936\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30805\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__30805\,
            I => \ADC_VDC.n22625\
        );

    \I__4934\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__30799\,
            I => \ADC_VDC.n6\
        );

    \I__4932\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30791\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__30795\,
            I => \N__30788\
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__30794\,
            I => \N__30785\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__30791\,
            I => \N__30782\
        );

    \I__4928\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30779\
        );

    \I__4927\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30776\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__30782\,
            I => \N__30773\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30768\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__30776\,
            I => \N__30768\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__30773\,
            I => cmd_rdadctmp_22_adj_1552
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__30768\,
            I => cmd_rdadctmp_22_adj_1552
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__30763\,
            I => \ADC_VDC.n11183_cascade_\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__30760\,
            I => \N__30757\
        );

    \I__4919\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30754\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__30754\,
            I => \N__30750\
        );

    \I__4917\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30747\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__30750\,
            I => \N__30744\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__30747\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__30744\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__4913\ : CEMux
    port map (
            O => \N__30739\,
            I => \N__30736\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__30736\,
            I => \N__30733\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__30733\,
            I => \N__30730\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__30730\,
            I => \N__30727\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__30727\,
            I => \ADC_VDC.n13957\
        );

    \I__4908\ : SRMux
    port map (
            O => \N__30724\,
            I => \N__30721\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30718\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__30718\,
            I => \ADC_VDC.n21707\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__30715\,
            I => \ADC_VDC.n17_cascade_\
        );

    \I__4904\ : InMux
    port map (
            O => \N__30712\,
            I => \N__30709\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__30709\,
            I => \N__30706\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__30706\,
            I => \ADC_VDC.n22055\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__30703\,
            I => \ADC_VDC.n27_cascade_\
        );

    \I__4900\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30697\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__30697\,
            I => \ADC_VDC.n10\
        );

    \I__4898\ : CEMux
    port map (
            O => \N__30694\,
            I => \N__30691\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__30691\,
            I => \N__30688\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__30688\,
            I => \ADC_VDC.n21869\
        );

    \I__4895\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30682\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__30682\,
            I => \ADC_VDC.n11923\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__30679\,
            I => \ADC_VDC.n11923_cascade_\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__30676\,
            I => \ADC_VDC.n20869_cascade_\
        );

    \I__4891\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__30670\,
            I => \N__30667\
        );

    \I__4889\ : Span4Mux_h
    port map (
            O => \N__30667\,
            I => \N__30664\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__30664\,
            I => \ADC_VDC.n8031\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__30661\,
            I => \N__30658\
        );

    \I__4886\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30655\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30652\
        );

    \I__4884\ : Odrv12
    port map (
            O => \N__30652\,
            I => \ADC_VDC.n23531\
        );

    \I__4883\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__30646\,
            I => \ADC_VDC.n20869\
        );

    \I__4881\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30640\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__30640\,
            I => \N__30635\
        );

    \I__4879\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30632\
        );

    \I__4878\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30629\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__30635\,
            I => \N__30626\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__30632\,
            I => buf_dds1_10
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__30629\,
            I => buf_dds1_10
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__30626\,
            I => buf_dds1_10
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__30619\,
            I => \N__30616\
        );

    \I__4872\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30613\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__30613\,
            I => n22160
        );

    \I__4870\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30607\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__30607\,
            I => \N__30604\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__30604\,
            I => \N__30600\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__30603\,
            I => \N__30596\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__30600\,
            I => \N__30593\
        );

    \I__4865\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30590\
        );

    \I__4864\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30587\
        );

    \I__4863\ : Sp12to4
    port map (
            O => \N__30593\,
            I => \N__30584\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__30590\,
            I => \N__30581\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__30587\,
            I => buf_adcdata_iac_18
        );

    \I__4860\ : Odrv12
    port map (
            O => \N__30584\,
            I => buf_adcdata_iac_18
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__30581\,
            I => buf_adcdata_iac_18
        );

    \I__4858\ : IoInMux
    port map (
            O => \N__30574\,
            I => \N__30571\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30568\
        );

    \I__4856\ : Span4Mux_s2_v
    port map (
            O => \N__30568\,
            I => \N__30565\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__30565\,
            I => \N__30561\
        );

    \I__4854\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30557\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__30561\,
            I => \N__30554\
        );

    \I__4852\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30551\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__30557\,
            I => \N__30548\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__30554\,
            I => \IAC_FLT0\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__30551\,
            I => \IAC_FLT0\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__30548\,
            I => \IAC_FLT0\
        );

    \I__4847\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30538\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__30538\,
            I => n22161
        );

    \I__4845\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30532\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30528\
        );

    \I__4843\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30525\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__30528\,
            I => \ADC_VDC.adc_state_3_N_1316_1\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__30525\,
            I => \ADC_VDC.adc_state_3_N_1316_1\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__30520\,
            I => \ADC_VDC.n22404_cascade_\
        );

    \I__4839\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30514\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__30514\,
            I => \ADC_VDC.n17\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__30511\,
            I => \N__30507\
        );

    \I__4836\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30503\
        );

    \I__4835\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30500\
        );

    \I__4834\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30497\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__30503\,
            I => cmd_rdadctmp_24
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__30500\,
            I => cmd_rdadctmp_24
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__30497\,
            I => cmd_rdadctmp_24
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__30490\,
            I => \N__30487\
        );

    \I__4829\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__30484\,
            I => \N__30481\
        );

    \I__4827\ : Span4Mux_h
    port map (
            O => \N__30481\,
            I => \N__30477\
        );

    \I__4826\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30474\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__30477\,
            I => cmd_rdadctmp_5
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__30474\,
            I => cmd_rdadctmp_5
        );

    \I__4823\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30466\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30463\
        );

    \I__4821\ : Odrv12
    port map (
            O => \N__30463\,
            I => n23468
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__4819\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30453\
        );

    \I__4818\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30449\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30446\
        );

    \I__4816\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30443\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__30449\,
            I => cmd_rdadctmp_25
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__30446\,
            I => cmd_rdadctmp_25
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__30443\,
            I => cmd_rdadctmp_25
        );

    \I__4812\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30429\
        );

    \I__4811\ : InMux
    port map (
            O => \N__30435\,
            I => \N__30426\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__30434\,
            I => \N__30419\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__30433\,
            I => \N__30415\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__30432\,
            I => \N__30412\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__30429\,
            I => \N__30405\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__30426\,
            I => \N__30405\
        );

    \I__4805\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30402\
        );

    \I__4804\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30395\
        );

    \I__4803\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30395\
        );

    \I__4802\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30395\
        );

    \I__4801\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30382\
        );

    \I__4800\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30382\
        );

    \I__4799\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30382\
        );

    \I__4798\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30382\
        );

    \I__4797\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30382\
        );

    \I__4796\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30382\
        );

    \I__4795\ : Odrv12
    port map (
            O => \N__30405\,
            I => \DTRIG_N_1182\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__30402\,
            I => \DTRIG_N_1182\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__30395\,
            I => \DTRIG_N_1182\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__30382\,
            I => \DTRIG_N_1182\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__30373\,
            I => \N__30368\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__30372\,
            I => \N__30362\
        );

    \I__4789\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30359\
        );

    \I__4788\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30356\
        );

    \I__4787\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30353\
        );

    \I__4786\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30346\
        );

    \I__4785\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30346\
        );

    \I__4784\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30346\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__30359\,
            I => \N__30337\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__30356\,
            I => \N__30334\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30331\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30328\
        );

    \I__4779\ : InMux
    port map (
            O => \N__30345\,
            I => \N__30315\
        );

    \I__4778\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30315\
        );

    \I__4777\ : InMux
    port map (
            O => \N__30343\,
            I => \N__30315\
        );

    \I__4776\ : InMux
    port map (
            O => \N__30342\,
            I => \N__30315\
        );

    \I__4775\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30315\
        );

    \I__4774\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30315\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__30337\,
            I => adc_state_1
        );

    \I__4772\ : Odrv12
    port map (
            O => \N__30334\,
            I => adc_state_1
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__30331\,
            I => adc_state_1
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__30328\,
            I => adc_state_1
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__30315\,
            I => adc_state_1
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__30304\,
            I => \N__30300\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__30303\,
            I => \N__30297\
        );

    \I__4766\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30294\
        );

    \I__4765\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30291\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30288\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30284\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30281\
        );

    \I__4761\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30278\
        );

    \I__4760\ : Odrv12
    port map (
            O => \N__30284\,
            I => cmd_rdadctmp_27
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__30281\,
            I => cmd_rdadctmp_27
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__30278\,
            I => cmd_rdadctmp_27
        );

    \I__4757\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30264\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__30267\,
            I => \N__30260\
        );

    \I__4754\ : Span12Mux_v
    port map (
            O => \N__30264\,
            I => \N__30257\
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__30263\,
            I => \N__30254\
        );

    \I__4752\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30251\
        );

    \I__4751\ : Span12Mux_h
    port map (
            O => \N__30257\,
            I => \N__30248\
        );

    \I__4750\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30245\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__30251\,
            I => buf_adcdata_iac_17
        );

    \I__4748\ : Odrv12
    port map (
            O => \N__30248\,
            I => buf_adcdata_iac_17
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__30245\,
            I => buf_adcdata_iac_17
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__30238\,
            I => \N__30235\
        );

    \I__4745\ : CascadeBuf
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__30232\,
            I => \N__30229\
        );

    \I__4743\ : CascadeBuf
    port map (
            O => \N__30229\,
            I => \N__30226\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__4741\ : CascadeBuf
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__4739\ : CascadeBuf
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \N__30211\
        );

    \I__4737\ : CascadeBuf
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__30208\,
            I => \N__30205\
        );

    \I__4735\ : CascadeBuf
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__30202\,
            I => \N__30199\
        );

    \I__4733\ : CascadeBuf
    port map (
            O => \N__30199\,
            I => \N__30196\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__4731\ : CascadeBuf
    port map (
            O => \N__30193\,
            I => \N__30190\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__30190\,
            I => \N__30186\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__30189\,
            I => \N__30183\
        );

    \I__4728\ : CascadeBuf
    port map (
            O => \N__30186\,
            I => \N__30180\
        );

    \I__4727\ : CascadeBuf
    port map (
            O => \N__30183\,
            I => \N__30177\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__30180\,
            I => \N__30174\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__30177\,
            I => \N__30171\
        );

    \I__4724\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30168\
        );

    \I__4723\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30165\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__30168\,
            I => \N__30162\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__30165\,
            I => \N__30158\
        );

    \I__4720\ : Span12Mux_s7_h
    port map (
            O => \N__30162\,
            I => \N__30155\
        );

    \I__4719\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30152\
        );

    \I__4718\ : Span12Mux_h
    port map (
            O => \N__30158\,
            I => \N__30147\
        );

    \I__4717\ : Span12Mux_h
    port map (
            O => \N__30155\,
            I => \N__30147\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30152\,
            I => data_count_6
        );

    \I__4715\ : Odrv12
    port map (
            O => \N__30147\,
            I => data_count_6
        );

    \I__4714\ : InMux
    port map (
            O => \N__30142\,
            I => n20618
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__30139\,
            I => \N__30136\
        );

    \I__4712\ : CascadeBuf
    port map (
            O => \N__30136\,
            I => \N__30133\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__4710\ : CascadeBuf
    port map (
            O => \N__30130\,
            I => \N__30127\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__30127\,
            I => \N__30124\
        );

    \I__4708\ : CascadeBuf
    port map (
            O => \N__30124\,
            I => \N__30121\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__30121\,
            I => \N__30118\
        );

    \I__4706\ : CascadeBuf
    port map (
            O => \N__30118\,
            I => \N__30115\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__30115\,
            I => \N__30112\
        );

    \I__4704\ : CascadeBuf
    port map (
            O => \N__30112\,
            I => \N__30109\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__30109\,
            I => \N__30106\
        );

    \I__4702\ : CascadeBuf
    port map (
            O => \N__30106\,
            I => \N__30103\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__30103\,
            I => \N__30100\
        );

    \I__4700\ : CascadeBuf
    port map (
            O => \N__30100\,
            I => \N__30097\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__30097\,
            I => \N__30094\
        );

    \I__4698\ : CascadeBuf
    port map (
            O => \N__30094\,
            I => \N__30090\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__30093\,
            I => \N__30087\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__30090\,
            I => \N__30084\
        );

    \I__4695\ : CascadeBuf
    port map (
            O => \N__30087\,
            I => \N__30081\
        );

    \I__4694\ : CascadeBuf
    port map (
            O => \N__30084\,
            I => \N__30078\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__30081\,
            I => \N__30075\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__30078\,
            I => \N__30072\
        );

    \I__4691\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30069\
        );

    \I__4690\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30066\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30063\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30060\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__30063\,
            I => \N__30057\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__30060\,
            I => \N__30054\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__30057\,
            I => \N__30050\
        );

    \I__4684\ : Sp12to4
    port map (
            O => \N__30054\,
            I => \N__30047\
        );

    \I__4683\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30044\
        );

    \I__4682\ : Sp12to4
    port map (
            O => \N__30050\,
            I => \N__30039\
        );

    \I__4681\ : Span12Mux_h
    port map (
            O => \N__30047\,
            I => \N__30039\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__30044\,
            I => data_count_7
        );

    \I__4679\ : Odrv12
    port map (
            O => \N__30039\,
            I => data_count_7
        );

    \I__4678\ : InMux
    port map (
            O => \N__30034\,
            I => n20619
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__30031\,
            I => \N__30028\
        );

    \I__4676\ : CascadeBuf
    port map (
            O => \N__30028\,
            I => \N__30025\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__30025\,
            I => \N__30022\
        );

    \I__4674\ : CascadeBuf
    port map (
            O => \N__30022\,
            I => \N__30019\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__30019\,
            I => \N__30016\
        );

    \I__4672\ : CascadeBuf
    port map (
            O => \N__30016\,
            I => \N__30013\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__30013\,
            I => \N__30010\
        );

    \I__4670\ : CascadeBuf
    port map (
            O => \N__30010\,
            I => \N__30007\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__30007\,
            I => \N__30004\
        );

    \I__4668\ : CascadeBuf
    port map (
            O => \N__30004\,
            I => \N__30001\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__4666\ : CascadeBuf
    port map (
            O => \N__29998\,
            I => \N__29995\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__29995\,
            I => \N__29992\
        );

    \I__4664\ : CascadeBuf
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__4662\ : CascadeBuf
    port map (
            O => \N__29986\,
            I => \N__29982\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__29985\,
            I => \N__29979\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__29982\,
            I => \N__29976\
        );

    \I__4659\ : CascadeBuf
    port map (
            O => \N__29979\,
            I => \N__29973\
        );

    \I__4658\ : CascadeBuf
    port map (
            O => \N__29976\,
            I => \N__29970\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__29973\,
            I => \N__29967\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__29970\,
            I => \N__29964\
        );

    \I__4655\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29961\
        );

    \I__4654\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29958\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__29961\,
            I => \N__29955\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29952\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__29955\,
            I => \N__29948\
        );

    \I__4650\ : Span12Mux_v
    port map (
            O => \N__29952\,
            I => \N__29945\
        );

    \I__4649\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29942\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__29948\,
            I => \N__29939\
        );

    \I__4647\ : Span12Mux_h
    port map (
            O => \N__29945\,
            I => \N__29936\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__29942\,
            I => data_count_8
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__29939\,
            I => data_count_8
        );

    \I__4644\ : Odrv12
    port map (
            O => \N__29936\,
            I => data_count_8
        );

    \I__4643\ : InMux
    port map (
            O => \N__29929\,
            I => \bfn_9_15_0_\
        );

    \I__4642\ : InMux
    port map (
            O => \N__29926\,
            I => n20621
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__29923\,
            I => \N__29920\
        );

    \I__4640\ : CascadeBuf
    port map (
            O => \N__29920\,
            I => \N__29917\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__29917\,
            I => \N__29914\
        );

    \I__4638\ : CascadeBuf
    port map (
            O => \N__29914\,
            I => \N__29911\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__29911\,
            I => \N__29908\
        );

    \I__4636\ : CascadeBuf
    port map (
            O => \N__29908\,
            I => \N__29905\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__29905\,
            I => \N__29902\
        );

    \I__4634\ : CascadeBuf
    port map (
            O => \N__29902\,
            I => \N__29899\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__29899\,
            I => \N__29896\
        );

    \I__4632\ : CascadeBuf
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__29893\,
            I => \N__29890\
        );

    \I__4630\ : CascadeBuf
    port map (
            O => \N__29890\,
            I => \N__29887\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__4628\ : CascadeBuf
    port map (
            O => \N__29884\,
            I => \N__29881\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__29881\,
            I => \N__29878\
        );

    \I__4626\ : CascadeBuf
    port map (
            O => \N__29878\,
            I => \N__29875\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__29875\,
            I => \N__29871\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__29874\,
            I => \N__29868\
        );

    \I__4623\ : CascadeBuf
    port map (
            O => \N__29871\,
            I => \N__29865\
        );

    \I__4622\ : CascadeBuf
    port map (
            O => \N__29868\,
            I => \N__29862\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__29865\,
            I => \N__29859\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__29862\,
            I => \N__29856\
        );

    \I__4619\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29853\
        );

    \I__4618\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29850\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29847\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__29850\,
            I => \N__29843\
        );

    \I__4615\ : Span12Mux_v
    port map (
            O => \N__29847\,
            I => \N__29840\
        );

    \I__4614\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29837\
        );

    \I__4613\ : Span12Mux_v
    port map (
            O => \N__29843\,
            I => \N__29834\
        );

    \I__4612\ : Span12Mux_h
    port map (
            O => \N__29840\,
            I => \N__29831\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__29837\,
            I => data_count_9
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__29834\,
            I => data_count_9
        );

    \I__4609\ : Odrv12
    port map (
            O => \N__29831\,
            I => data_count_9
        );

    \I__4608\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29821\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__29821\,
            I => \N__29818\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__29818\,
            I => n11983
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__29815\,
            I => \n24_adj_1598_cascade_\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__29812\,
            I => \n24_adj_1506_cascade_\
        );

    \I__4603\ : IoInMux
    port map (
            O => \N__29809\,
            I => \N__29806\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29803\
        );

    \I__4601\ : Span4Mux_s2_v
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__4600\ : Span4Mux_h
    port map (
            O => \N__29800\,
            I => \N__29796\
        );

    \I__4599\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29793\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__29796\,
            I => \N__29790\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29786\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__29790\,
            I => \N__29783\
        );

    \I__4595\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29780\
        );

    \I__4594\ : Span4Mux_h
    port map (
            O => \N__29786\,
            I => \N__29777\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__29783\,
            I => \IAC_FLT1\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__29780\,
            I => \IAC_FLT1\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__29777\,
            I => \IAC_FLT1\
        );

    \I__4590\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29767\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__29767\,
            I => n11982
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__29764\,
            I => \N__29761\
        );

    \I__4587\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29758\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__29758\,
            I => \N__29754\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__29757\,
            I => \N__29751\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__29754\,
            I => \N__29747\
        );

    \I__4583\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29744\
        );

    \I__4582\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29741\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__29747\,
            I => cmd_rdadctmp_18
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__29744\,
            I => cmd_rdadctmp_18
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__29741\,
            I => cmd_rdadctmp_18
        );

    \I__4578\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29729\
        );

    \I__4577\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29726\
        );

    \I__4576\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29723\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29720\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29717\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__29723\,
            I => buf_dds1_11
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__29720\,
            I => buf_dds1_11
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__29717\,
            I => buf_dds1_11
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__29710\,
            I => \N__29707\
        );

    \I__4569\ : CascadeBuf
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__29704\,
            I => \N__29701\
        );

    \I__4567\ : CascadeBuf
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__29698\,
            I => \N__29695\
        );

    \I__4565\ : CascadeBuf
    port map (
            O => \N__29695\,
            I => \N__29692\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__29692\,
            I => \N__29689\
        );

    \I__4563\ : CascadeBuf
    port map (
            O => \N__29689\,
            I => \N__29686\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__4561\ : CascadeBuf
    port map (
            O => \N__29683\,
            I => \N__29680\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__4559\ : CascadeBuf
    port map (
            O => \N__29677\,
            I => \N__29674\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29671\
        );

    \I__4557\ : CascadeBuf
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__29668\,
            I => \N__29665\
        );

    \I__4555\ : CascadeBuf
    port map (
            O => \N__29665\,
            I => \N__29661\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__29664\,
            I => \N__29658\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__29661\,
            I => \N__29655\
        );

    \I__4552\ : CascadeBuf
    port map (
            O => \N__29658\,
            I => \N__29652\
        );

    \I__4551\ : CascadeBuf
    port map (
            O => \N__29655\,
            I => \N__29649\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__29652\,
            I => \N__29646\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__29649\,
            I => \N__29643\
        );

    \I__4548\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29640\
        );

    \I__4547\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29637\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29634\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29631\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__29634\,
            I => \N__29627\
        );

    \I__4543\ : Span12Mux_v
    port map (
            O => \N__29631\,
            I => \N__29624\
        );

    \I__4542\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29621\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__29627\,
            I => \N__29618\
        );

    \I__4540\ : Span12Mux_h
    port map (
            O => \N__29624\,
            I => \N__29615\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__29621\,
            I => data_count_0
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__29618\,
            I => data_count_0
        );

    \I__4537\ : Odrv12
    port map (
            O => \N__29615\,
            I => data_count_0
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__29608\,
            I => \N__29605\
        );

    \I__4535\ : CascadeBuf
    port map (
            O => \N__29605\,
            I => \N__29602\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__29602\,
            I => \N__29599\
        );

    \I__4533\ : CascadeBuf
    port map (
            O => \N__29599\,
            I => \N__29596\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__29596\,
            I => \N__29593\
        );

    \I__4531\ : CascadeBuf
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__29590\,
            I => \N__29587\
        );

    \I__4529\ : CascadeBuf
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__4527\ : CascadeBuf
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__4526\ : CascadeMux
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__4525\ : CascadeBuf
    port map (
            O => \N__29575\,
            I => \N__29572\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__29572\,
            I => \N__29569\
        );

    \I__4523\ : CascadeBuf
    port map (
            O => \N__29569\,
            I => \N__29566\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__29566\,
            I => \N__29563\
        );

    \I__4521\ : CascadeBuf
    port map (
            O => \N__29563\,
            I => \N__29560\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__29560\,
            I => \N__29557\
        );

    \I__4519\ : CascadeBuf
    port map (
            O => \N__29557\,
            I => \N__29553\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__29556\,
            I => \N__29550\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__29553\,
            I => \N__29547\
        );

    \I__4516\ : CascadeBuf
    port map (
            O => \N__29550\,
            I => \N__29544\
        );

    \I__4515\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29541\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__29544\,
            I => \N__29538\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29535\
        );

    \I__4512\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29532\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__29535\,
            I => \N__29529\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__29532\,
            I => \N__29526\
        );

    \I__4509\ : Span4Mux_h
    port map (
            O => \N__29529\,
            I => \N__29523\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__29526\,
            I => \N__29519\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__29523\,
            I => \N__29516\
        );

    \I__4506\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29513\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__29519\,
            I => \N__29510\
        );

    \I__4504\ : Span4Mux_h
    port map (
            O => \N__29516\,
            I => \N__29507\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__29513\,
            I => data_count_1
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__29510\,
            I => data_count_1
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__29507\,
            I => data_count_1
        );

    \I__4500\ : InMux
    port map (
            O => \N__29500\,
            I => n20613
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__29497\,
            I => \N__29494\
        );

    \I__4498\ : CascadeBuf
    port map (
            O => \N__29494\,
            I => \N__29491\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__29491\,
            I => \N__29488\
        );

    \I__4496\ : CascadeBuf
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__29485\,
            I => \N__29482\
        );

    \I__4494\ : CascadeBuf
    port map (
            O => \N__29482\,
            I => \N__29479\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__29479\,
            I => \N__29476\
        );

    \I__4492\ : CascadeBuf
    port map (
            O => \N__29476\,
            I => \N__29473\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \N__29470\
        );

    \I__4490\ : CascadeBuf
    port map (
            O => \N__29470\,
            I => \N__29467\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__29467\,
            I => \N__29464\
        );

    \I__4488\ : CascadeBuf
    port map (
            O => \N__29464\,
            I => \N__29461\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__4486\ : CascadeBuf
    port map (
            O => \N__29458\,
            I => \N__29455\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__4484\ : CascadeBuf
    port map (
            O => \N__29452\,
            I => \N__29449\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__29449\,
            I => \N__29445\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__29448\,
            I => \N__29442\
        );

    \I__4481\ : CascadeBuf
    port map (
            O => \N__29445\,
            I => \N__29439\
        );

    \I__4480\ : CascadeBuf
    port map (
            O => \N__29442\,
            I => \N__29436\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__29439\,
            I => \N__29433\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \N__29430\
        );

    \I__4477\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29427\
        );

    \I__4476\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29424\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29421\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__29424\,
            I => \N__29418\
        );

    \I__4473\ : Sp12to4
    port map (
            O => \N__29421\,
            I => \N__29415\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__29418\,
            I => \N__29411\
        );

    \I__4471\ : Span12Mux_v
    port map (
            O => \N__29415\,
            I => \N__29408\
        );

    \I__4470\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29405\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__29411\,
            I => \N__29402\
        );

    \I__4468\ : Span12Mux_h
    port map (
            O => \N__29408\,
            I => \N__29399\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__29405\,
            I => data_count_2
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__29402\,
            I => data_count_2
        );

    \I__4465\ : Odrv12
    port map (
            O => \N__29399\,
            I => data_count_2
        );

    \I__4464\ : InMux
    port map (
            O => \N__29392\,
            I => n20614
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__29389\,
            I => \N__29386\
        );

    \I__4462\ : CascadeBuf
    port map (
            O => \N__29386\,
            I => \N__29383\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__29383\,
            I => \N__29380\
        );

    \I__4460\ : CascadeBuf
    port map (
            O => \N__29380\,
            I => \N__29377\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__4458\ : CascadeBuf
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__4456\ : CascadeBuf
    port map (
            O => \N__29368\,
            I => \N__29365\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__29365\,
            I => \N__29362\
        );

    \I__4454\ : CascadeBuf
    port map (
            O => \N__29362\,
            I => \N__29359\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__29359\,
            I => \N__29356\
        );

    \I__4452\ : CascadeBuf
    port map (
            O => \N__29356\,
            I => \N__29353\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__29353\,
            I => \N__29350\
        );

    \I__4450\ : CascadeBuf
    port map (
            O => \N__29350\,
            I => \N__29347\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \N__29344\
        );

    \I__4448\ : CascadeBuf
    port map (
            O => \N__29344\,
            I => \N__29340\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__29343\,
            I => \N__29337\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__29340\,
            I => \N__29334\
        );

    \I__4445\ : CascadeBuf
    port map (
            O => \N__29337\,
            I => \N__29331\
        );

    \I__4444\ : CascadeBuf
    port map (
            O => \N__29334\,
            I => \N__29328\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__29331\,
            I => \N__29325\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__29328\,
            I => \N__29322\
        );

    \I__4441\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29319\
        );

    \I__4440\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29316\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29313\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29310\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__29313\,
            I => \N__29306\
        );

    \I__4436\ : Span12Mux_v
    port map (
            O => \N__29310\,
            I => \N__29303\
        );

    \I__4435\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29300\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__29306\,
            I => \N__29297\
        );

    \I__4433\ : Span12Mux_h
    port map (
            O => \N__29303\,
            I => \N__29294\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__29300\,
            I => data_count_3
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__29297\,
            I => data_count_3
        );

    \I__4430\ : Odrv12
    port map (
            O => \N__29294\,
            I => data_count_3
        );

    \I__4429\ : InMux
    port map (
            O => \N__29287\,
            I => n20615
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__29284\,
            I => \N__29281\
        );

    \I__4427\ : CascadeBuf
    port map (
            O => \N__29281\,
            I => \N__29278\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__29278\,
            I => \N__29275\
        );

    \I__4425\ : CascadeBuf
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__29272\,
            I => \N__29269\
        );

    \I__4423\ : CascadeBuf
    port map (
            O => \N__29269\,
            I => \N__29266\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__4421\ : CascadeBuf
    port map (
            O => \N__29263\,
            I => \N__29260\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \N__29257\
        );

    \I__4419\ : CascadeBuf
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__29254\,
            I => \N__29251\
        );

    \I__4417\ : CascadeBuf
    port map (
            O => \N__29251\,
            I => \N__29248\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__29248\,
            I => \N__29245\
        );

    \I__4415\ : CascadeBuf
    port map (
            O => \N__29245\,
            I => \N__29242\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__29242\,
            I => \N__29239\
        );

    \I__4413\ : CascadeBuf
    port map (
            O => \N__29239\,
            I => \N__29235\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__29238\,
            I => \N__29232\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__29235\,
            I => \N__29229\
        );

    \I__4410\ : CascadeBuf
    port map (
            O => \N__29232\,
            I => \N__29226\
        );

    \I__4409\ : CascadeBuf
    port map (
            O => \N__29229\,
            I => \N__29223\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__29226\,
            I => \N__29220\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__29223\,
            I => \N__29217\
        );

    \I__4406\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29214\
        );

    \I__4405\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29211\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__29211\,
            I => \N__29205\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__29208\,
            I => \N__29202\
        );

    \I__4401\ : Sp12to4
    port map (
            O => \N__29205\,
            I => \N__29199\
        );

    \I__4400\ : Span4Mux_h
    port map (
            O => \N__29202\,
            I => \N__29195\
        );

    \I__4399\ : Span12Mux_s8_v
    port map (
            O => \N__29199\,
            I => \N__29192\
        );

    \I__4398\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29189\
        );

    \I__4397\ : Sp12to4
    port map (
            O => \N__29195\,
            I => \N__29184\
        );

    \I__4396\ : Span12Mux_h
    port map (
            O => \N__29192\,
            I => \N__29184\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__29189\,
            I => data_count_4
        );

    \I__4394\ : Odrv12
    port map (
            O => \N__29184\,
            I => data_count_4
        );

    \I__4393\ : InMux
    port map (
            O => \N__29179\,
            I => n20616
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__29176\,
            I => \N__29173\
        );

    \I__4391\ : CascadeBuf
    port map (
            O => \N__29173\,
            I => \N__29170\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__29170\,
            I => \N__29167\
        );

    \I__4389\ : CascadeBuf
    port map (
            O => \N__29167\,
            I => \N__29164\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__29164\,
            I => \N__29161\
        );

    \I__4387\ : CascadeBuf
    port map (
            O => \N__29161\,
            I => \N__29158\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__29158\,
            I => \N__29155\
        );

    \I__4385\ : CascadeBuf
    port map (
            O => \N__29155\,
            I => \N__29152\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__29152\,
            I => \N__29149\
        );

    \I__4383\ : CascadeBuf
    port map (
            O => \N__29149\,
            I => \N__29146\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__29146\,
            I => \N__29143\
        );

    \I__4381\ : CascadeBuf
    port map (
            O => \N__29143\,
            I => \N__29140\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__29140\,
            I => \N__29137\
        );

    \I__4379\ : CascadeBuf
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__29134\,
            I => \N__29131\
        );

    \I__4377\ : CascadeBuf
    port map (
            O => \N__29131\,
            I => \N__29127\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__29130\,
            I => \N__29124\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__29127\,
            I => \N__29121\
        );

    \I__4374\ : CascadeBuf
    port map (
            O => \N__29124\,
            I => \N__29118\
        );

    \I__4373\ : CascadeBuf
    port map (
            O => \N__29121\,
            I => \N__29115\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29112\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__29115\,
            I => \N__29109\
        );

    \I__4370\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29106\
        );

    \I__4369\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29103\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__29106\,
            I => \N__29100\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29097\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__29100\,
            I => \N__29093\
        );

    \I__4365\ : Span12Mux_s7_v
    port map (
            O => \N__29097\,
            I => \N__29090\
        );

    \I__4364\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29087\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__29093\,
            I => \N__29084\
        );

    \I__4362\ : Span12Mux_h
    port map (
            O => \N__29090\,
            I => \N__29081\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__29087\,
            I => data_count_5
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__29084\,
            I => data_count_5
        );

    \I__4359\ : Odrv12
    port map (
            O => \N__29081\,
            I => data_count_5
        );

    \I__4358\ : InMux
    port map (
            O => \N__29074\,
            I => n20617
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__29071\,
            I => \n22164_cascade_\
        );

    \I__4356\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29063\
        );

    \I__4355\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29060\
        );

    \I__4354\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29057\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29054\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__29060\,
            I => buf_dds1_14
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__29057\,
            I => buf_dds1_14
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__29054\,
            I => buf_dds1_14
        );

    \I__4349\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29044\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__29044\,
            I => \N__29041\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__29041\,
            I => \N__29038\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__29038\,
            I => n23366
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__29035\,
            I => \n16_adj_1763_cascade_\
        );

    \I__4344\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29029\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__29029\,
            I => n23369
        );

    \I__4342\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29023\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__29023\,
            I => \N__29020\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__29020\,
            I => \N__29017\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__29017\,
            I => \N__29014\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__29014\,
            I => n30_adj_1698
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__29011\,
            I => \N__29005\
        );

    \I__4336\ : InMux
    port map (
            O => \N__29010\,
            I => \N__28998\
        );

    \I__4335\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28998\
        );

    \I__4334\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28998\
        );

    \I__4333\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28995\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__28998\,
            I => \N__28991\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__28995\,
            I => \N__28988\
        );

    \I__4330\ : CascadeMux
    port map (
            O => \N__28994\,
            I => \N__28985\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28982\
        );

    \I__4328\ : Span12Mux_h
    port map (
            O => \N__28988\,
            I => \N__28979\
        );

    \I__4327\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28976\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__28982\,
            I => \N__28973\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__28979\,
            I => \buf_cfgRTD_6\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__28976\,
            I => \buf_cfgRTD_6\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__28973\,
            I => \buf_cfgRTD_6\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__28966\,
            I => \N__28962\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__28965\,
            I => \N__28959\
        );

    \I__4320\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28954\
        );

    \I__4319\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28954\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28950\
        );

    \I__4317\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28947\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__28950\,
            I => \N__28942\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__28947\,
            I => \N__28942\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__28942\,
            I => \N__28937\
        );

    \I__4313\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28934\
        );

    \I__4312\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28931\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__28937\,
            I => \buf_cfgRTD_2\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__28934\,
            I => \buf_cfgRTD_2\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__28931\,
            I => \buf_cfgRTD_2\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__28924\,
            I => \N__28919\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__28923\,
            I => \N__28916\
        );

    \I__4306\ : InMux
    port map (
            O => \N__28922\,
            I => \N__28911\
        );

    \I__4305\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28911\
        );

    \I__4304\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28908\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28905\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__28908\,
            I => \N__28902\
        );

    \I__4301\ : Span4Mux_v
    port map (
            O => \N__28905\,
            I => \N__28895\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__28902\,
            I => \N__28895\
        );

    \I__4299\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28892\
        );

    \I__4298\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28889\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__28895\,
            I => \N__28884\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__28892\,
            I => \N__28884\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__28889\,
            I => \buf_cfgRTD_4\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__28884\,
            I => \buf_cfgRTD_4\
        );

    \I__4293\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28876\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__28876\,
            I => \N__28872\
        );

    \I__4291\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28869\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__28872\,
            I => \comm_spi.n24028\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__28869\,
            I => \comm_spi.n24028\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__28864\,
            I => \comm_spi.n24028_cascade_\
        );

    \I__4287\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__4284\ : Span4Mux_v
    port map (
            O => \N__28852\,
            I => \N__28848\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__28851\,
            I => \N__28845\
        );

    \I__4282\ : Sp12to4
    port map (
            O => \N__28848\,
            I => \N__28842\
        );

    \I__4281\ : InMux
    port map (
            O => \N__28845\,
            I => \N__28839\
        );

    \I__4280\ : Odrv12
    port map (
            O => \N__28842\,
            I => \buf_readRTD_12\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__28839\,
            I => \buf_readRTD_12\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__28834\,
            I => \N__28831\
        );

    \I__4277\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28828\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__28828\,
            I => n20_adj_1781
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__28825\,
            I => \N__28822\
        );

    \I__4274\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28818\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__28821\,
            I => \N__28815\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28812\
        );

    \I__4271\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28809\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__28812\,
            I => \N__28806\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28802\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__28806\,
            I => \N__28799\
        );

    \I__4267\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28796\
        );

    \I__4266\ : Odrv12
    port map (
            O => \N__28802\,
            I => cmd_rdadctmp_19_adj_1529
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__28799\,
            I => cmd_rdadctmp_19_adj_1529
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__28796\,
            I => cmd_rdadctmp_19_adj_1529
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28785\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__28788\,
            I => \N__28782\
        );

    \I__4261\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28779\
        );

    \I__4260\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28776\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__28779\,
            I => \N__28773\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__28776\,
            I => \N__28770\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__28773\,
            I => \N__28764\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__28770\,
            I => \N__28764\
        );

    \I__4255\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28761\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__28764\,
            I => cmd_rdadctmp_20_adj_1528
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__28761\,
            I => cmd_rdadctmp_20_adj_1528
        );

    \I__4252\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28753\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__28753\,
            I => n23309
        );

    \I__4250\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__4247\ : Sp12to4
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__28740\,
            I => \N__28734\
        );

    \I__4245\ : Span12Mux_h
    port map (
            O => \N__28737\,
            I => \N__28731\
        );

    \I__4244\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28728\
        );

    \I__4243\ : Odrv12
    port map (
            O => \N__28731\,
            I => \buf_readRTD_10\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__28728\,
            I => \buf_readRTD_10\
        );

    \I__4241\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28719\
        );

    \I__4240\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28715\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__28719\,
            I => \N__28712\
        );

    \I__4238\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28709\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__28715\,
            I => \N__28706\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__28712\,
            I => \N__28703\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__28709\,
            I => buf_dds1_5
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__28706\,
            I => buf_dds1_5
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__28703\,
            I => buf_dds1_5
        );

    \I__4232\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__28693\,
            I => \N__28689\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__28692\,
            I => \N__28686\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__28689\,
            I => \N__28683\
        );

    \I__4228\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28680\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__28683\,
            I => buf_adcdata_vdc_14
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__28680\,
            I => buf_adcdata_vdc_14
        );

    \I__4225\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28672\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28668\
        );

    \I__4223\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28665\
        );

    \I__4222\ : Span12Mux_s10_h
    port map (
            O => \N__28668\,
            I => \N__28661\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__28665\,
            I => \N__28658\
        );

    \I__4220\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28655\
        );

    \I__4219\ : Span12Mux_h
    port map (
            O => \N__28661\,
            I => \N__28652\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__28658\,
            I => \N__28649\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__28655\,
            I => buf_adcdata_vac_14
        );

    \I__4216\ : Odrv12
    port map (
            O => \N__28652\,
            I => buf_adcdata_vac_14
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__28649\,
            I => buf_adcdata_vac_14
        );

    \I__4214\ : CEMux
    port map (
            O => \N__28642\,
            I => \N__28639\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__28639\,
            I => \N__28633\
        );

    \I__4212\ : CEMux
    port map (
            O => \N__28638\,
            I => \N__28630\
        );

    \I__4211\ : CEMux
    port map (
            O => \N__28637\,
            I => \N__28627\
        );

    \I__4210\ : CEMux
    port map (
            O => \N__28636\,
            I => \N__28622\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__28633\,
            I => \N__28616\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28616\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__28627\,
            I => \N__28613\
        );

    \I__4206\ : CEMux
    port map (
            O => \N__28626\,
            I => \N__28610\
        );

    \I__4205\ : CEMux
    port map (
            O => \N__28625\,
            I => \N__28607\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__28622\,
            I => \N__28604\
        );

    \I__4203\ : CEMux
    port map (
            O => \N__28621\,
            I => \N__28601\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__28616\,
            I => \N__28598\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__28613\,
            I => \N__28593\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__28610\,
            I => \N__28593\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__28607\,
            I => \N__28590\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__28604\,
            I => \N__28582\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28582\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__28598\,
            I => \N__28582\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__28593\,
            I => \N__28579\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__28590\,
            I => \N__28576\
        );

    \I__4193\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28573\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__28582\,
            I => \ADC_VDC.n14120\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__28579\,
            I => \ADC_VDC.n14120\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__28576\,
            I => \ADC_VDC.n14120\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__28573\,
            I => \ADC_VDC.n14120\
        );

    \I__4188\ : SRMux
    port map (
            O => \N__28564\,
            I => \N__28558\
        );

    \I__4187\ : SRMux
    port map (
            O => \N__28563\,
            I => \N__28554\
        );

    \I__4186\ : SRMux
    port map (
            O => \N__28562\,
            I => \N__28550\
        );

    \I__4185\ : SRMux
    port map (
            O => \N__28561\,
            I => \N__28546\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__28558\,
            I => \N__28543\
        );

    \I__4183\ : SRMux
    port map (
            O => \N__28557\,
            I => \N__28540\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28537\
        );

    \I__4181\ : SRMux
    port map (
            O => \N__28553\,
            I => \N__28534\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__28550\,
            I => \N__28531\
        );

    \I__4179\ : SRMux
    port map (
            O => \N__28549\,
            I => \N__28528\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28525\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__28543\,
            I => \N__28522\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__28540\,
            I => \N__28519\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__28537\,
            I => \N__28516\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28513\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__28531\,
            I => \N__28510\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__28528\,
            I => \N__28507\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__28525\,
            I => \N__28504\
        );

    \I__4170\ : Span4Mux_v
    port map (
            O => \N__28522\,
            I => \N__28497\
        );

    \I__4169\ : Span4Mux_h
    port map (
            O => \N__28519\,
            I => \N__28497\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__28516\,
            I => \N__28497\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__28513\,
            I => \N__28492\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__28510\,
            I => \N__28492\
        );

    \I__4165\ : Odrv12
    port map (
            O => \N__28507\,
            I => \ADC_VDC.n15721\
        );

    \I__4164\ : Odrv4
    port map (
            O => \N__28504\,
            I => \ADC_VDC.n15721\
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__28497\,
            I => \ADC_VDC.n15721\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__28492\,
            I => \ADC_VDC.n15721\
        );

    \I__4161\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__28480\,
            I => \ADC_VDC.cmd_rdadcbuf_35_N_1344_34\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__28477\,
            I => \ADC_VDC.n4_cascade_\
        );

    \I__4158\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__28468\,
            I => \N__28463\
        );

    \I__4155\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28460\
        );

    \I__4154\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28457\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__28463\,
            I => cmd_rdadcbuf_34
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__28460\,
            I => cmd_rdadcbuf_34
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__28457\,
            I => cmd_rdadcbuf_34
        );

    \I__4150\ : CEMux
    port map (
            O => \N__28450\,
            I => \N__28447\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28444\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__28444\,
            I => \N__28441\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__28441\,
            I => \ADC_VDC.n14092\
        );

    \I__4146\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28434\
        );

    \I__4145\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28431\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__28434\,
            I => cmd_rdadcbuf_14
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__28431\,
            I => cmd_rdadcbuf_14
        );

    \I__4142\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28422\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__28425\,
            I => \N__28418\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__28422\,
            I => \N__28415\
        );

    \I__4139\ : InMux
    port map (
            O => \N__28421\,
            I => \N__28412\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28409\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__28415\,
            I => cmd_rdadctmp_8_adj_1566
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__28412\,
            I => cmd_rdadctmp_8_adj_1566
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__28409\,
            I => cmd_rdadctmp_8_adj_1566
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__28402\,
            I => \N__28398\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__28401\,
            I => \N__28387\
        );

    \I__4132\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28382\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__28397\,
            I => \N__28376\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__28396\,
            I => \N__28373\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \N__28367\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__28394\,
            I => \N__28364\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__28393\,
            I => \N__28361\
        );

    \I__4126\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28348\
        );

    \I__4125\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28348\
        );

    \I__4124\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28348\
        );

    \I__4123\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28348\
        );

    \I__4122\ : InMux
    port map (
            O => \N__28386\,
            I => \N__28348\
        );

    \I__4121\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28348\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__28382\,
            I => \N__28345\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__28381\,
            I => \N__28339\
        );

    \I__4118\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28328\
        );

    \I__4117\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28328\
        );

    \I__4116\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28328\
        );

    \I__4115\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28328\
        );

    \I__4114\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28315\
        );

    \I__4113\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28315\
        );

    \I__4112\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28315\
        );

    \I__4111\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28315\
        );

    \I__4110\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28315\
        );

    \I__4109\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28315\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__28348\,
            I => \N__28310\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__28345\,
            I => \N__28310\
        );

    \I__4106\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28297\
        );

    \I__4105\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28297\
        );

    \I__4104\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28297\
        );

    \I__4103\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28297\
        );

    \I__4102\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28297\
        );

    \I__4101\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28297\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__28328\,
            I => \N__28292\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__28315\,
            I => \N__28292\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__28310\,
            I => n13925
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__28297\,
            I => n13925
        );

    \I__4096\ : Odrv12
    port map (
            O => \N__28292\,
            I => n13925
        );

    \I__4095\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28278\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__28281\,
            I => \N__28274\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__28278\,
            I => \N__28271\
        );

    \I__4091\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28268\
        );

    \I__4090\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28265\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__28271\,
            I => cmd_rdadctmp_9_adj_1565
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__28268\,
            I => cmd_rdadctmp_9_adj_1565
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__28265\,
            I => cmd_rdadctmp_9_adj_1565
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__28258\,
            I => \N__28255\
        );

    \I__4085\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28251\
        );

    \I__4084\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28248\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__28251\,
            I => cmd_rdadcbuf_22
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__28248\,
            I => cmd_rdadcbuf_22
        );

    \I__4081\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28239\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28236\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28239\,
            I => cmd_rdadcbuf_13
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__28236\,
            I => cmd_rdadcbuf_13
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__4076\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28224\
        );

    \I__4075\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28221\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__28224\,
            I => cmd_rdadcbuf_16
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__28221\,
            I => cmd_rdadcbuf_16
        );

    \I__4072\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__28207\,
            I => \N__28203\
        );

    \I__4068\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28200\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__28203\,
            I => buf_adcdata_vdc_5
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__28200\,
            I => buf_adcdata_vdc_5
        );

    \I__4065\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28188\
        );

    \I__4063\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28185\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__28188\,
            I => cmd_rdadcbuf_27
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__28185\,
            I => cmd_rdadcbuf_27
        );

    \I__4060\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28176\
        );

    \I__4059\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__28176\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__28173\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4056\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28165\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__28165\,
            I => \N__28162\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__28162\,
            I => \ADC_VDC.n20\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__28159\,
            I => \ADC_VDC.n19_cascade_\
        );

    \I__4052\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__28150\,
            I => \ADC_VDC.n21\
        );

    \I__4049\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28144\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__28144\,
            I => \ADC_VDC.n28\
        );

    \I__4047\ : CEMux
    port map (
            O => \N__28141\,
            I => \N__28138\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__28135\,
            I => \ADC_VDC.n21871\
        );

    \I__4044\ : CEMux
    port map (
            O => \N__28132\,
            I => \N__28129\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__28129\,
            I => \ADC_VDC.n13865\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__28126\,
            I => \ADC_VDC.n9_cascade_\
        );

    \I__4041\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28118\
        );

    \I__4040\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28113\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28113\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__28118\,
            I => \ADC_VDC.n22071\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__28113\,
            I => \ADC_VDC.n22071\
        );

    \I__4036\ : SRMux
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28102\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__28102\,
            I => \N__28099\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__28099\,
            I => \ADC_VDC.n5\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__28096\,
            I => \N__28093\
        );

    \I__4031\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28085\
        );

    \I__4029\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28080\
        );

    \I__4028\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28080\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__28085\,
            I => cmd_rdadctmp_21
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__28080\,
            I => cmd_rdadctmp_21
        );

    \I__4025\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28070\
        );

    \I__4024\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28065\
        );

    \I__4023\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28065\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__28070\,
            I => cmd_rdadctmp_22
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__28065\,
            I => cmd_rdadctmp_22
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__28060\,
            I => \N__28056\
        );

    \I__4019\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28048\
        );

    \I__4018\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28048\
        );

    \I__4017\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28048\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__28048\,
            I => cmd_rdadctmp_23
        );

    \I__4015\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28041\
        );

    \I__4014\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28038\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__28041\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__28038\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__4011\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28029\
        );

    \I__4010\ : InMux
    port map (
            O => \N__28032\,
            I => \N__28026\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__28029\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__28026\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__4006\ : InMux
    port map (
            O => \N__28018\,
            I => \N__28014\
        );

    \I__4005\ : InMux
    port map (
            O => \N__28017\,
            I => \N__28011\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__28014\,
            I => \N__28008\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__28011\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__28008\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__4001\ : InMux
    port map (
            O => \N__28003\,
            I => \N__28000\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__27994\,
            I => \N__27989\
        );

    \I__3997\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27986\
        );

    \I__3996\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27983\
        );

    \I__3995\ : Sp12to4
    port map (
            O => \N__27989\,
            I => \N__27980\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27977\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__27983\,
            I => buf_adcdata_iac_19
        );

    \I__3992\ : Odrv12
    port map (
            O => \N__27980\,
            I => buf_adcdata_iac_19
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__27977\,
            I => buf_adcdata_iac_19
        );

    \I__3990\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27965\
        );

    \I__3989\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27962\
        );

    \I__3988\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27959\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27956\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__27962\,
            I => \N__27953\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__27959\,
            I => buf_dds1_12
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__27956\,
            I => buf_dds1_12
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__27953\,
            I => buf_dds1_12
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__27946\,
            I => \N__27943\
        );

    \I__3981\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27940\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__3979\ : Odrv4
    port map (
            O => \N__27937\,
            I => n16_adj_1778
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__27934\,
            I => \N__27931\
        );

    \I__3977\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27928\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__27928\,
            I => \N__27923\
        );

    \I__3975\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27918\
        );

    \I__3974\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27918\
        );

    \I__3973\ : Odrv12
    port map (
            O => \N__27923\,
            I => cmd_rdadctmp_26
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__27918\,
            I => cmd_rdadctmp_26
        );

    \I__3971\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27910\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__27910\,
            I => \N__27905\
        );

    \I__3969\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27902\
        );

    \I__3968\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27899\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__27905\,
            I => \N__27896\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__27902\,
            I => buf_dds1_7
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__27899\,
            I => buf_dds1_7
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__27896\,
            I => buf_dds1_7
        );

    \I__3963\ : IoInMux
    port map (
            O => \N__27889\,
            I => \N__27886\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27882\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__3960\ : Span12Mux_s9_v
    port map (
            O => \N__27882\,
            I => \N__27876\
        );

    \I__3959\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27873\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__27876\,
            I => \IAC_SCLK\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__27873\,
            I => \IAC_SCLK\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__3955\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__27862\,
            I => \N__27858\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__27861\,
            I => \N__27855\
        );

    \I__3952\ : Span4Mux_v
    port map (
            O => \N__27858\,
            I => \N__27851\
        );

    \I__3951\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27846\
        );

    \I__3950\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27846\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__27851\,
            I => cmd_rdadctmp_27_adj_1521
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__27846\,
            I => cmd_rdadctmp_27_adj_1521
        );

    \I__3947\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__27829\,
            I => \N__27825\
        );

    \I__3942\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27821\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__27825\,
            I => \N__27818\
        );

    \I__3940\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27815\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__27821\,
            I => buf_adcdata_vac_19
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__27818\,
            I => buf_adcdata_vac_19
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__27815\,
            I => buf_adcdata_vac_19
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__27808\,
            I => \n23474_cascade_\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__27805\,
            I => \n23477_cascade_\
        );

    \I__3934\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27799\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__27799\,
            I => n30_adj_1784
        );

    \I__3932\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27793\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27790\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__27790\,
            I => n112_adj_1772
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__27787\,
            I => \n30_adj_1768_cascade_\
        );

    \I__3928\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27781\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__27781\,
            I => n19_adj_1780
        );

    \I__3926\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27775\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__27775\,
            I => \N__27772\
        );

    \I__3924\ : Span4Mux_h
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__3923\ : Span4Mux_h
    port map (
            O => \N__27769\,
            I => \N__27766\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__27766\,
            I => n30_adj_1702
        );

    \I__3921\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27760\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__27760\,
            I => n22358
        );

    \I__3919\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27754\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__27754\,
            I => \N__27750\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__27753\,
            I => \N__27747\
        );

    \I__3916\ : Span4Mux_v
    port map (
            O => \N__27750\,
            I => \N__27744\
        );

    \I__3915\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27741\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__27744\,
            I => buf_adcdata_vdc_19
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__27741\,
            I => buf_adcdata_vdc_19
        );

    \I__3912\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27733\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__27733\,
            I => n19_adj_1789
        );

    \I__3910\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__27727\,
            I => n23426
        );

    \I__3908\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27721\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__27721\,
            I => n23429
        );

    \I__3906\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27714\
        );

    \I__3905\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27711\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__27714\,
            I => cmd_rdadcbuf_28
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__27711\,
            I => cmd_rdadcbuf_28
        );

    \I__3902\ : InMux
    port map (
            O => \N__27706\,
            I => \ADC_VDC.n20717\
        );

    \I__3901\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27699\
        );

    \I__3900\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27696\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__27699\,
            I => cmd_rdadcbuf_29
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__27696\,
            I => cmd_rdadcbuf_29
        );

    \I__3897\ : InMux
    port map (
            O => \N__27691\,
            I => \ADC_VDC.n20718\
        );

    \I__3896\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27684\
        );

    \I__3895\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27681\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__27684\,
            I => cmd_rdadcbuf_30
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__27681\,
            I => cmd_rdadcbuf_30
        );

    \I__3892\ : InMux
    port map (
            O => \N__27676\,
            I => \ADC_VDC.n20719\
        );

    \I__3891\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27669\
        );

    \I__3890\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27666\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__27669\,
            I => cmd_rdadcbuf_31
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__27666\,
            I => cmd_rdadcbuf_31
        );

    \I__3887\ : InMux
    port map (
            O => \N__27661\,
            I => \ADC_VDC.n20720\
        );

    \I__3886\ : InMux
    port map (
            O => \N__27658\,
            I => \bfn_8_10_0_\
        );

    \I__3885\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27651\
        );

    \I__3884\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27648\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__27651\,
            I => cmd_rdadcbuf_33
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__27648\,
            I => cmd_rdadcbuf_33
        );

    \I__3881\ : InMux
    port map (
            O => \N__27643\,
            I => \ADC_VDC.n20722\
        );

    \I__3880\ : InMux
    port map (
            O => \N__27640\,
            I => \ADC_VDC.n20723\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__27637\,
            I => \N__27632\
        );

    \I__3878\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27627\
        );

    \I__3877\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27627\
        );

    \I__3876\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27624\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__27627\,
            I => cmd_rdadctmp_20_adj_1554
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__27624\,
            I => cmd_rdadctmp_20_adj_1554
        );

    \I__3873\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27616\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27612\
        );

    \I__3871\ : InMux
    port map (
            O => \N__27615\,
            I => \N__27609\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__27612\,
            I => cmd_rdadcbuf_20
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__27609\,
            I => cmd_rdadcbuf_20
        );

    \I__3868\ : InMux
    port map (
            O => \N__27604\,
            I => \ADC_VDC.n20709\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__27601\,
            I => \N__27596\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__27600\,
            I => \N__27593\
        );

    \I__3865\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27590\
        );

    \I__3864\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27587\
        );

    \I__3863\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27584\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__27590\,
            I => cmd_rdadctmp_21_adj_1553
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__27587\,
            I => cmd_rdadctmp_21_adj_1553
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__27584\,
            I => cmd_rdadctmp_21_adj_1553
        );

    \I__3859\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27573\
        );

    \I__3858\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27570\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__27573\,
            I => \N__27567\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27564\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__27567\,
            I => cmd_rdadcbuf_21
        );

    \I__3854\ : Odrv4
    port map (
            O => \N__27564\,
            I => cmd_rdadcbuf_21
        );

    \I__3853\ : InMux
    port map (
            O => \N__27559\,
            I => \ADC_VDC.n20710\
        );

    \I__3852\ : InMux
    port map (
            O => \N__27556\,
            I => \ADC_VDC.n20711\
        );

    \I__3851\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27549\
        );

    \I__3850\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27546\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__27549\,
            I => cmd_rdadcbuf_23
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__27546\,
            I => cmd_rdadcbuf_23
        );

    \I__3847\ : InMux
    port map (
            O => \N__27541\,
            I => \ADC_VDC.n20712\
        );

    \I__3846\ : InMux
    port map (
            O => \N__27538\,
            I => \bfn_8_9_0_\
        );

    \I__3845\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27531\
        );

    \I__3844\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27528\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__27531\,
            I => cmd_rdadcbuf_25
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__27528\,
            I => cmd_rdadcbuf_25
        );

    \I__3841\ : InMux
    port map (
            O => \N__27523\,
            I => \ADC_VDC.n20714\
        );

    \I__3840\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27516\
        );

    \I__3839\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27513\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__27516\,
            I => cmd_rdadcbuf_26
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__27513\,
            I => cmd_rdadcbuf_26
        );

    \I__3836\ : InMux
    port map (
            O => \N__27508\,
            I => \ADC_VDC.n20715\
        );

    \I__3835\ : InMux
    port map (
            O => \N__27505\,
            I => \ADC_VDC.n20716\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__27502\,
            I => \N__27497\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__27501\,
            I => \N__27494\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__27500\,
            I => \N__27491\
        );

    \I__3831\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27488\
        );

    \I__3830\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27485\
        );

    \I__3829\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27482\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__27488\,
            I => cmd_rdadctmp_12_adj_1562
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__27485\,
            I => cmd_rdadctmp_12_adj_1562
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__27482\,
            I => cmd_rdadctmp_12_adj_1562
        );

    \I__3825\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27471\
        );

    \I__3824\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27468\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__27471\,
            I => cmd_rdadcbuf_12
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__27468\,
            I => cmd_rdadcbuf_12
        );

    \I__3821\ : InMux
    port map (
            O => \N__27463\,
            I => \ADC_VDC.n20701\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \N__27455\
        );

    \I__3819\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27450\
        );

    \I__3818\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27450\
        );

    \I__3817\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27447\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__27450\,
            I => cmd_rdadctmp_13_adj_1561
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__27447\,
            I => cmd_rdadctmp_13_adj_1561
        );

    \I__3814\ : InMux
    port map (
            O => \N__27442\,
            I => \ADC_VDC.n20702\
        );

    \I__3813\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27434\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27431\
        );

    \I__3811\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27428\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__27434\,
            I => \N__27425\
        );

    \I__3809\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27422\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__27428\,
            I => cmd_rdadctmp_14_adj_1560
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__27425\,
            I => cmd_rdadctmp_14_adj_1560
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__27422\,
            I => cmd_rdadctmp_14_adj_1560
        );

    \I__3805\ : InMux
    port map (
            O => \N__27415\,
            I => \ADC_VDC.n20703\
        );

    \I__3804\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27407\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__27411\,
            I => \N__27404\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__27410\,
            I => \N__27401\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27398\
        );

    \I__3800\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27395\
        );

    \I__3799\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27392\
        );

    \I__3798\ : Span4Mux_v
    port map (
            O => \N__27398\,
            I => \N__27389\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27386\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__27392\,
            I => cmd_rdadctmp_15_adj_1559
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__27389\,
            I => cmd_rdadctmp_15_adj_1559
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__27386\,
            I => cmd_rdadctmp_15_adj_1559
        );

    \I__3793\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27376\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__27376\,
            I => \N__27372\
        );

    \I__3791\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27369\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__27372\,
            I => cmd_rdadcbuf_15
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__27369\,
            I => cmd_rdadcbuf_15
        );

    \I__3788\ : InMux
    port map (
            O => \N__27364\,
            I => \ADC_VDC.n20704\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__27361\,
            I => \N__27356\
        );

    \I__3786\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27353\
        );

    \I__3785\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27350\
        );

    \I__3784\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27347\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__27353\,
            I => cmd_rdadctmp_16_adj_1558
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__27350\,
            I => cmd_rdadctmp_16_adj_1558
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__27347\,
            I => cmd_rdadctmp_16_adj_1558
        );

    \I__3780\ : InMux
    port map (
            O => \N__27340\,
            I => \bfn_8_8_0_\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__27337\,
            I => \N__27333\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__27336\,
            I => \N__27329\
        );

    \I__3777\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27326\
        );

    \I__3776\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27323\
        );

    \I__3775\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27320\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__27326\,
            I => cmd_rdadctmp_17_adj_1557
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__27323\,
            I => cmd_rdadctmp_17_adj_1557
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__27320\,
            I => cmd_rdadctmp_17_adj_1557
        );

    \I__3771\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27310\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27306\
        );

    \I__3769\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27303\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__27306\,
            I => cmd_rdadcbuf_17
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__27303\,
            I => cmd_rdadcbuf_17
        );

    \I__3766\ : InMux
    port map (
            O => \N__27298\,
            I => \ADC_VDC.n20706\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__27295\,
            I => \N__27290\
        );

    \I__3764\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27285\
        );

    \I__3763\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27285\
        );

    \I__3762\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27282\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__27285\,
            I => cmd_rdadctmp_18_adj_1556
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__27282\,
            I => cmd_rdadctmp_18_adj_1556
        );

    \I__3759\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27273\
        );

    \I__3758\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27270\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__27273\,
            I => cmd_rdadcbuf_18
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__27270\,
            I => cmd_rdadcbuf_18
        );

    \I__3755\ : InMux
    port map (
            O => \N__27265\,
            I => \ADC_VDC.n20707\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__27262\,
            I => \N__27257\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__27261\,
            I => \N__27254\
        );

    \I__3752\ : InMux
    port map (
            O => \N__27260\,
            I => \N__27251\
        );

    \I__3751\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27248\
        );

    \I__3750\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27245\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__27251\,
            I => cmd_rdadctmp_19_adj_1555
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__27248\,
            I => cmd_rdadctmp_19_adj_1555
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27245\,
            I => cmd_rdadctmp_19_adj_1555
        );

    \I__3746\ : InMux
    port map (
            O => \N__27238\,
            I => \N__27235\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27231\
        );

    \I__3744\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27228\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__27231\,
            I => cmd_rdadcbuf_19
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27228\,
            I => cmd_rdadcbuf_19
        );

    \I__3741\ : InMux
    port map (
            O => \N__27223\,
            I => \ADC_VDC.n20708\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__27220\,
            I => \N__27215\
        );

    \I__3739\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27210\
        );

    \I__3738\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27210\
        );

    \I__3737\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27207\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__27210\,
            I => cmd_rdadctmp_4_adj_1570
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__27207\,
            I => cmd_rdadctmp_4_adj_1570
        );

    \I__3734\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27199\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__27199\,
            I => \ADC_VDC.cmd_rdadcbuf_4\
        );

    \I__3732\ : InMux
    port map (
            O => \N__27196\,
            I => \ADC_VDC.n20693\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__27193\,
            I => \N__27189\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__27192\,
            I => \N__27185\
        );

    \I__3729\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27180\
        );

    \I__3728\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27180\
        );

    \I__3727\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27177\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__27180\,
            I => cmd_rdadctmp_5_adj_1569
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__27177\,
            I => cmd_rdadctmp_5_adj_1569
        );

    \I__3724\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__27169\,
            I => \N__27166\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__27166\,
            I => \ADC_VDC.cmd_rdadcbuf_5\
        );

    \I__3721\ : InMux
    port map (
            O => \N__27163\,
            I => \ADC_VDC.n20694\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__27160\,
            I => \N__27155\
        );

    \I__3719\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27152\
        );

    \I__3718\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27149\
        );

    \I__3717\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27146\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__27152\,
            I => cmd_rdadctmp_6_adj_1568
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27149\,
            I => cmd_rdadctmp_6_adj_1568
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__27146\,
            I => cmd_rdadctmp_6_adj_1568
        );

    \I__3713\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__27136\,
            I => \ADC_VDC.cmd_rdadcbuf_6\
        );

    \I__3711\ : InMux
    port map (
            O => \N__27133\,
            I => \ADC_VDC.n20695\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__27130\,
            I => \N__27125\
        );

    \I__3709\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27120\
        );

    \I__3708\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27120\
        );

    \I__3707\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27117\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__27120\,
            I => cmd_rdadctmp_7_adj_1567
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__27117\,
            I => cmd_rdadctmp_7_adj_1567
        );

    \I__3704\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__27109\,
            I => \ADC_VDC.cmd_rdadcbuf_7\
        );

    \I__3702\ : InMux
    port map (
            O => \N__27106\,
            I => \ADC_VDC.n20696\
        );

    \I__3701\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27100\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__27100\,
            I => \ADC_VDC.cmd_rdadcbuf_8\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27097\,
            I => \bfn_8_7_0_\
        );

    \I__3698\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27091\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__27091\,
            I => \ADC_VDC.cmd_rdadcbuf_9\
        );

    \I__3696\ : InMux
    port map (
            O => \N__27088\,
            I => \ADC_VDC.n20698\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__27085\,
            I => \N__27080\
        );

    \I__3694\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27077\
        );

    \I__3693\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27074\
        );

    \I__3692\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27071\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__27077\,
            I => cmd_rdadctmp_10_adj_1564
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__27074\,
            I => cmd_rdadctmp_10_adj_1564
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__27071\,
            I => cmd_rdadctmp_10_adj_1564
        );

    \I__3688\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__27061\,
            I => \ADC_VDC.cmd_rdadcbuf_10\
        );

    \I__3686\ : InMux
    port map (
            O => \N__27058\,
            I => \ADC_VDC.n20699\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__27055\,
            I => \N__27050\
        );

    \I__3684\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27045\
        );

    \I__3683\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27045\
        );

    \I__3682\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27042\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__27045\,
            I => cmd_rdadctmp_11_adj_1563
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__27042\,
            I => cmd_rdadctmp_11_adj_1563
        );

    \I__3679\ : InMux
    port map (
            O => \N__27037\,
            I => \ADC_VDC.n20700\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__27034\,
            I => \N__27029\
        );

    \I__3677\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27026\
        );

    \I__3676\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27023\
        );

    \I__3675\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27020\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__27026\,
            I => cmd_rdadctmp_0_adj_1574
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__27023\,
            I => cmd_rdadctmp_0_adj_1574
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__27020\,
            I => cmd_rdadctmp_0_adj_1574
        );

    \I__3671\ : InMux
    port map (
            O => \N__27013\,
            I => \N__27010\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__27010\,
            I => \ADC_VDC.cmd_rdadcbuf_0\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__27007\,
            I => \N__27002\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__27006\,
            I => \N__26999\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__27005\,
            I => \N__26996\
        );

    \I__3666\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26991\
        );

    \I__3665\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26991\
        );

    \I__3664\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26988\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__26991\,
            I => cmd_rdadctmp_1_adj_1573
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__26988\,
            I => cmd_rdadctmp_1_adj_1573
        );

    \I__3661\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26980\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__26980\,
            I => \ADC_VDC.cmd_rdadcbuf_1\
        );

    \I__3659\ : InMux
    port map (
            O => \N__26977\,
            I => \ADC_VDC.n20690\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__3657\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26966\
        );

    \I__3656\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26963\
        );

    \I__3655\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26960\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26957\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__26963\,
            I => cmd_rdadctmp_2_adj_1572
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__26960\,
            I => cmd_rdadctmp_2_adj_1572
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__26957\,
            I => cmd_rdadctmp_2_adj_1572
        );

    \I__3650\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26947\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__26947\,
            I => \ADC_VDC.cmd_rdadcbuf_2\
        );

    \I__3648\ : InMux
    port map (
            O => \N__26944\,
            I => \ADC_VDC.n20691\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \N__26936\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__26940\,
            I => \N__26933\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__26939\,
            I => \N__26930\
        );

    \I__3644\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26925\
        );

    \I__3643\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26925\
        );

    \I__3642\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26922\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__26925\,
            I => cmd_rdadctmp_3_adj_1571
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__26922\,
            I => cmd_rdadctmp_3_adj_1571
        );

    \I__3639\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26914\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__26914\,
            I => \ADC_VDC.cmd_rdadcbuf_3\
        );

    \I__3637\ : InMux
    port map (
            O => \N__26911\,
            I => \ADC_VDC.n20692\
        );

    \I__3636\ : InMux
    port map (
            O => \N__26908\,
            I => \bfn_8_3_0_\
        );

    \I__3635\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26901\
        );

    \I__3634\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26898\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__26901\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__26898\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__3631\ : InMux
    port map (
            O => \N__26893\,
            I => \ADC_VDC.n20733\
        );

    \I__3630\ : InMux
    port map (
            O => \N__26890\,
            I => \ADC_VDC.n20734\
        );

    \I__3629\ : InMux
    port map (
            O => \N__26887\,
            I => \ADC_VDC.n20735\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__26884\,
            I => \N__26881\
        );

    \I__3627\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26877\
        );

    \I__3626\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26874\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26871\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__26874\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__26871\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__3622\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26859\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__26865\,
            I => \N__26849\
        );

    \I__3620\ : InMux
    port map (
            O => \N__26864\,
            I => \N__26843\
        );

    \I__3619\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26840\
        );

    \I__3618\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26834\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__26859\,
            I => \N__26831\
        );

    \I__3616\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26828\
        );

    \I__3615\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26823\
        );

    \I__3614\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26823\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__26855\,
            I => \N__26819\
        );

    \I__3612\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26814\
        );

    \I__3611\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26805\
        );

    \I__3610\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26805\
        );

    \I__3609\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26805\
        );

    \I__3608\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26805\
        );

    \I__3607\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26800\
        );

    \I__3606\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26800\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__26843\,
            I => \N__26795\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26792\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__26839\,
            I => \N__26787\
        );

    \I__3602\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26782\
        );

    \I__3601\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26779\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26772\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__26831\,
            I => \N__26772\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26772\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26768\
        );

    \I__3596\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26765\
        );

    \I__3595\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26762\
        );

    \I__3594\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26759\
        );

    \I__3593\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26756\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__26814\,
            I => \N__26749\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26749\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26749\
        );

    \I__3589\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26746\
        );

    \I__3588\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26743\
        );

    \I__3587\ : Span4Mux_h
    port map (
            O => \N__26795\,
            I => \N__26738\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__26792\,
            I => \N__26738\
        );

    \I__3585\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26733\
        );

    \I__3584\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26733\
        );

    \I__3583\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26726\
        );

    \I__3582\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26726\
        );

    \I__3581\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26726\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__26782\,
            I => \N__26721\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__26779\,
            I => \N__26721\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__26772\,
            I => \N__26718\
        );

    \I__3577\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26715\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__26768\,
            I => \N__26710\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26710\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__26762\,
            I => \N__26701\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__26759\,
            I => \N__26701\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__26756\,
            I => \N__26701\
        );

    \I__3571\ : Span12Mux_h
    port map (
            O => \N__26749\,
            I => \N__26701\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__26746\,
            I => \RTD.adc_state_3\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__26743\,
            I => \RTD.adc_state_3\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__26738\,
            I => \RTD.adc_state_3\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__26733\,
            I => \RTD.adc_state_3\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__26726\,
            I => \RTD.adc_state_3\
        );

    \I__3565\ : Odrv12
    port map (
            O => \N__26721\,
            I => \RTD.adc_state_3\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__26718\,
            I => \RTD.adc_state_3\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__26715\,
            I => \RTD.adc_state_3\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__26710\,
            I => \RTD.adc_state_3\
        );

    \I__3561\ : Odrv12
    port map (
            O => \N__26701\,
            I => \RTD.adc_state_3\
        );

    \I__3560\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26664\
        );

    \I__3558\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26661\
        );

    \I__3557\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26658\
        );

    \I__3556\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26655\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__26673\,
            I => \N__26647\
        );

    \I__3554\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26643\
        );

    \I__3553\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26632\
        );

    \I__3552\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26632\
        );

    \I__3551\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26632\
        );

    \I__3550\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26632\
        );

    \I__3549\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26632\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__26664\,
            I => \N__26625\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N__26625\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26625\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__26655\,
            I => \N__26622\
        );

    \I__3544\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26619\
        );

    \I__3543\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26613\
        );

    \I__3542\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26610\
        );

    \I__3541\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26599\
        );

    \I__3540\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26599\
        );

    \I__3539\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26594\
        );

    \I__3538\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26594\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26591\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__26632\,
            I => \N__26588\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__26625\,
            I => \N__26581\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__26622\,
            I => \N__26581\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__26619\,
            I => \N__26581\
        );

    \I__3532\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26574\
        );

    \I__3531\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26574\
        );

    \I__3530\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26574\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26569\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26569\
        );

    \I__3527\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26566\
        );

    \I__3526\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26561\
        );

    \I__3525\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26561\
        );

    \I__3524\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26556\
        );

    \I__3523\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26556\
        );

    \I__3522\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26553\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__26599\,
            I => \N__26550\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__26594\,
            I => \N__26547\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__26591\,
            I => \N__26536\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__26588\,
            I => \N__26536\
        );

    \I__3517\ : Span4Mux_h
    port map (
            O => \N__26581\,
            I => \N__26536\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__26574\,
            I => \N__26536\
        );

    \I__3515\ : Span4Mux_h
    port map (
            O => \N__26569\,
            I => \N__26536\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__26566\,
            I => \RTD.adc_state_1\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__26561\,
            I => \RTD.adc_state_1\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__26556\,
            I => \RTD.adc_state_1\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__26553\,
            I => \RTD.adc_state_1\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__26550\,
            I => \RTD.adc_state_1\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__26547\,
            I => \RTD.adc_state_1\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__26536\,
            I => \RTD.adc_state_1\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__26521\,
            I => \N__26511\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__26520\,
            I => \N__26507\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \N__26504\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__26518\,
            I => \N__26487\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__26517\,
            I => \N__26483\
        );

    \I__3502\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26476\
        );

    \I__3501\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26476\
        );

    \I__3500\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26476\
        );

    \I__3499\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26469\
        );

    \I__3498\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26466\
        );

    \I__3497\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26463\
        );

    \I__3496\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26460\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__26503\,
            I => \N__26456\
        );

    \I__3494\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26441\
        );

    \I__3493\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26441\
        );

    \I__3492\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26441\
        );

    \I__3491\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26441\
        );

    \I__3490\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26441\
        );

    \I__3489\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26441\
        );

    \I__3488\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26441\
        );

    \I__3487\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26438\
        );

    \I__3486\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26425\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26425\
        );

    \I__3484\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26418\
        );

    \I__3483\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26418\
        );

    \I__3482\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26418\
        );

    \I__3481\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26415\
        );

    \I__3480\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26412\
        );

    \I__3479\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26409\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__26476\,
            I => \N__26406\
        );

    \I__3477\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26399\
        );

    \I__3476\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26399\
        );

    \I__3475\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26399\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__26472\,
            I => \N__26395\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__26469\,
            I => \N__26389\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__26466\,
            I => \N__26382\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26382\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__26460\,
            I => \N__26382\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \N__26379\
        );

    \I__3468\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26376\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__26441\,
            I => \N__26367\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26367\
        );

    \I__3465\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26356\
        );

    \I__3464\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26356\
        );

    \I__3463\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26356\
        );

    \I__3462\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26356\
        );

    \I__3461\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26356\
        );

    \I__3460\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26349\
        );

    \I__3459\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26349\
        );

    \I__3458\ : InMux
    port map (
            O => \N__26430\,
            I => \N__26349\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__26425\,
            I => \N__26340\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__26418\,
            I => \N__26340\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26340\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__26412\,
            I => \N__26340\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26337\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__26406\,
            I => \N__26332\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26332\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__26398\,
            I => \N__26329\
        );

    \I__3449\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26326\
        );

    \I__3448\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26323\
        );

    \I__3447\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26318\
        );

    \I__3446\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26318\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__26389\,
            I => \N__26313\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__26382\,
            I => \N__26313\
        );

    \I__3443\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26310\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26307\
        );

    \I__3441\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26298\
        );

    \I__3440\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26298\
        );

    \I__3439\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26298\
        );

    \I__3438\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26298\
        );

    \I__3437\ : Span12Mux_h
    port map (
            O => \N__26367\,
            I => \N__26291\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26291\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__26349\,
            I => \N__26291\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__26340\,
            I => \N__26284\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__26337\,
            I => \N__26284\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__26332\,
            I => \N__26284\
        );

    \I__3431\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26281\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26278\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__26323\,
            I => adc_state_2
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__26318\,
            I => adc_state_2
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__26313\,
            I => adc_state_2
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__26310\,
            I => adc_state_2
        );

    \I__3425\ : Odrv12
    port map (
            O => \N__26307\,
            I => adc_state_2
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__26298\,
            I => adc_state_2
        );

    \I__3423\ : Odrv12
    port map (
            O => \N__26291\,
            I => adc_state_2
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__26284\,
            I => adc_state_2
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__26281\,
            I => adc_state_2
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__26278\,
            I => adc_state_2
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26239\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26239\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26239\
        );

    \I__3415\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26239\
        );

    \I__3414\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26236\
        );

    \I__3413\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26230\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__26248\,
            I => \N__26226\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26217\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__26236\,
            I => \N__26217\
        );

    \I__3409\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26214\
        );

    \I__3408\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26210\
        );

    \I__3407\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26207\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26203\
        );

    \I__3405\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26200\
        );

    \I__3404\ : InMux
    port map (
            O => \N__26226\,
            I => \N__26197\
        );

    \I__3403\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26194\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__26224\,
            I => \N__26182\
        );

    \I__3401\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26178\
        );

    \I__3400\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26175\
        );

    \I__3399\ : Span4Mux_h
    port map (
            O => \N__26217\,
            I => \N__26169\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26169\
        );

    \I__3397\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26166\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N__26160\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26160\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26157\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__26203\,
            I => \N__26152\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__26200\,
            I => \N__26152\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__26197\,
            I => \N__26147\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__26194\,
            I => \N__26147\
        );

    \I__3389\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26127\
        );

    \I__3388\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26127\
        );

    \I__3387\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26127\
        );

    \I__3386\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26127\
        );

    \I__3385\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26127\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26127\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26127\
        );

    \I__3382\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26127\
        );

    \I__3381\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26124\
        );

    \I__3380\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26121\
        );

    \I__3379\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26118\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26114\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__26175\,
            I => \N__26111\
        );

    \I__3376\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26108\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__26169\,
            I => \N__26103\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__26166\,
            I => \N__26103\
        );

    \I__3373\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26100\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__26160\,
            I => \N__26097\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26092\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__26152\,
            I => \N__26092\
        );

    \I__3369\ : Span4Mux_v
    port map (
            O => \N__26147\,
            I => \N__26089\
        );

    \I__3368\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26082\
        );

    \I__3367\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26082\
        );

    \I__3366\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26082\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26077\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__26124\,
            I => \N__26077\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26072\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__26118\,
            I => \N__26072\
        );

    \I__3361\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26069\
        );

    \I__3360\ : Span4Mux_h
    port map (
            O => \N__26114\,
            I => \N__26060\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__26111\,
            I => \N__26060\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26060\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__26103\,
            I => \N__26060\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__26100\,
            I => \RTD.adc_state_0\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__26097\,
            I => \RTD.adc_state_0\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__26092\,
            I => \RTD.adc_state_0\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__26089\,
            I => \RTD.adc_state_0\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__26082\,
            I => \RTD.adc_state_0\
        );

    \I__3351\ : Odrv12
    port map (
            O => \N__26077\,
            I => \RTD.adc_state_0\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__26072\,
            I => \RTD.adc_state_0\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26069\,
            I => \RTD.adc_state_0\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__26060\,
            I => \RTD.adc_state_0\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__26041\,
            I => \ADC_VDC.n22071_cascade_\
        );

    \I__3346\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__3344\ : Span12Mux_h
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__3343\ : Odrv12
    port map (
            O => \N__26029\,
            I => \EIS_SYNCCLK\
        );

    \I__3342\ : IoInMux
    port map (
            O => \N__26026\,
            I => \N__26022\
        );

    \I__3341\ : IoInMux
    port map (
            O => \N__26025\,
            I => \N__26019\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__26016\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__26019\,
            I => \N__26013\
        );

    \I__3338\ : Span4Mux_s3_h
    port map (
            O => \N__26016\,
            I => \N__26010\
        );

    \I__3337\ : Span4Mux_s3_v
    port map (
            O => \N__26013\,
            I => \N__26007\
        );

    \I__3336\ : Span4Mux_h
    port map (
            O => \N__26010\,
            I => \N__26004\
        );

    \I__3335\ : Span4Mux_h
    port map (
            O => \N__26007\,
            I => \N__26001\
        );

    \I__3334\ : Span4Mux_h
    port map (
            O => \N__26004\,
            I => \N__25998\
        );

    \I__3333\ : Sp12to4
    port map (
            O => \N__26001\,
            I => \N__25993\
        );

    \I__3332\ : Sp12to4
    port map (
            O => \N__25998\,
            I => \N__25993\
        );

    \I__3331\ : Span12Mux_v
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__3330\ : Odrv12
    port map (
            O => \N__25990\,
            I => \IAC_CLK\
        );

    \I__3329\ : InMux
    port map (
            O => \N__25987\,
            I => \bfn_8_2_0_\
        );

    \I__3328\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25980\
        );

    \I__3327\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25977\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__25980\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__25977\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__3324\ : InMux
    port map (
            O => \N__25972\,
            I => \ADC_VDC.n20725\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__25969\,
            I => \N__25965\
        );

    \I__3322\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25962\
        );

    \I__3321\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25959\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__25962\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__25959\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__3318\ : InMux
    port map (
            O => \N__25954\,
            I => \ADC_VDC.n20726\
        );

    \I__3317\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25947\
        );

    \I__3316\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25944\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__25947\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__25944\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__3313\ : InMux
    port map (
            O => \N__25939\,
            I => \ADC_VDC.n20727\
        );

    \I__3312\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25932\
        );

    \I__3311\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25929\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__25932\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__25929\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__3308\ : InMux
    port map (
            O => \N__25924\,
            I => \ADC_VDC.n20728\
        );

    \I__3307\ : InMux
    port map (
            O => \N__25921\,
            I => \ADC_VDC.n20729\
        );

    \I__3306\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25914\
        );

    \I__3305\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25911\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__25914\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__25911\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__3302\ : InMux
    port map (
            O => \N__25906\,
            I => \ADC_VDC.n20730\
        );

    \I__3301\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25899\
        );

    \I__3300\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25896\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__25899\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__25896\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3297\ : InMux
    port map (
            O => \N__25891\,
            I => \ADC_VDC.n20731\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__25888\,
            I => \ADC_IAC.n22384_cascade_\
        );

    \I__3295\ : CEMux
    port map (
            O => \N__25885\,
            I => \N__25882\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__25882\,
            I => \N__25879\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__25879\,
            I => \ADC_IAC.n22032\
        );

    \I__3292\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25870\
        );

    \I__3291\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25870\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__25870\,
            I => \N__25864\
        );

    \I__3289\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25859\
        );

    \I__3288\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25859\
        );

    \I__3287\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25856\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__25864\,
            I => \N__25853\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__25859\,
            I => \N__25850\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__25856\,
            I => acadc_trig
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__25853\,
            I => acadc_trig
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__25850\,
            I => acadc_trig
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__25843\,
            I => \ADC_IAC.n17_cascade_\
        );

    \I__3280\ : CEMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__25834\,
            I => \ADC_IAC.n12\
        );

    \I__3277\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__25828\,
            I => n21892
        );

    \I__3275\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25822\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__25822\,
            I => n14_adj_1578
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__25819\,
            I => \N__25813\
        );

    \I__3272\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25807\
        );

    \I__3271\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25807\
        );

    \I__3270\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25802\
        );

    \I__3269\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25802\
        );

    \I__3268\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25799\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__25807\,
            I => \N__25796\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25793\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25790\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__25796\,
            I => \N__25787\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__25793\,
            I => \N__25782\
        );

    \I__3262\ : Span4Mux_v
    port map (
            O => \N__25790\,
            I => \N__25782\
        );

    \I__3261\ : Sp12to4
    port map (
            O => \N__25787\,
            I => \N__25777\
        );

    \I__3260\ : Sp12to4
    port map (
            O => \N__25782\,
            I => \N__25777\
        );

    \I__3259\ : Span12Mux_h
    port map (
            O => \N__25777\,
            I => \N__25774\
        );

    \I__3258\ : Odrv12
    port map (
            O => \N__25774\,
            I => \IAC_DRDY\
        );

    \I__3257\ : IoInMux
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__3255\ : Span12Mux_s8_v
    port map (
            O => \N__25765\,
            I => \N__25761\
        );

    \I__3254\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25758\
        );

    \I__3253\ : Odrv12
    port map (
            O => \N__25761\,
            I => \IAC_CS\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__25758\,
            I => \IAC_CS\
        );

    \I__3251\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__3250\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25747\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__25747\,
            I => cmd_rdadctmp_2
        );

    \I__3248\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25738\
        );

    \I__3247\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25738\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__25738\,
            I => cmd_rdadctmp_3
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__25735\,
            I => \N__25731\
        );

    \I__3244\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25726\
        );

    \I__3243\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25726\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__25726\,
            I => cmd_rdadctmp_4
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__3240\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25716\
        );

    \I__3239\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25713\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__25716\,
            I => cmd_rdadctmp_0
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__25713\,
            I => cmd_rdadctmp_0
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__3235\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__3234\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25699\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__25699\,
            I => cmd_rdadctmp_1
        );

    \I__3232\ : InMux
    port map (
            O => \N__25696\,
            I => \ADC_IAC.n20680\
        );

    \I__3231\ : InMux
    port map (
            O => \N__25693\,
            I => \ADC_IAC.n20681\
        );

    \I__3230\ : InMux
    port map (
            O => \N__25690\,
            I => \ADC_IAC.n20682\
        );

    \I__3229\ : CEMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__25684\,
            I => \N__25681\
        );

    \I__3227\ : Span4Mux_v
    port map (
            O => \N__25681\,
            I => \N__25678\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__25678\,
            I => \N__25674\
        );

    \I__3225\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__25674\,
            I => \ADC_IAC.n13667\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__25671\,
            I => \ADC_IAC.n13667\
        );

    \I__3222\ : SRMux
    port map (
            O => \N__25666\,
            I => \N__25663\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__25657\,
            I => \ADC_IAC.n15622\
        );

    \I__3218\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25651\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__25651\,
            I => \ADC_IAC.n22031\
        );

    \I__3216\ : InMux
    port map (
            O => \N__25648\,
            I => \N__25644\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25641\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__25644\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__25641\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3212\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25632\
        );

    \I__3211\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25629\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__25632\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__25629\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__25624\,
            I => \N__25620\
        );

    \I__3207\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25617\
        );

    \I__3206\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25614\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__25617\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__25614\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3203\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25605\
        );

    \I__3202\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25602\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__25605\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25602\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3199\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25593\
        );

    \I__3198\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25590\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__25593\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__25590\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3195\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25581\
        );

    \I__3194\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25578\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__25581\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__25578\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__25573\,
            I => \ADC_IAC.n22113_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25566\
        );

    \I__3189\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25563\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__25566\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__25563\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3186\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25554\
        );

    \I__3185\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25551\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__25554\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__25551\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \ADC_IAC.n22128_cascade_\
        );

    \I__3181\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25540\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__25540\,
            I => \N__25537\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__25537\,
            I => n19
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__25534\,
            I => \N__25531\
        );

    \I__3177\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25528\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__3175\ : Span4Mux_v
    port map (
            O => \N__25525\,
            I => \N__25521\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__25524\,
            I => \N__25518\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__25521\,
            I => \N__25515\
        );

    \I__3172\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25512\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__25515\,
            I => \buf_readRTD_0\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__25512\,
            I => \buf_readRTD_0\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__25507\,
            I => \n22041_cascade_\
        );

    \I__3168\ : InMux
    port map (
            O => \N__25504\,
            I => \bfn_7_16_0_\
        );

    \I__3167\ : InMux
    port map (
            O => \N__25501\,
            I => \ADC_IAC.n20676\
        );

    \I__3166\ : InMux
    port map (
            O => \N__25498\,
            I => \ADC_IAC.n20677\
        );

    \I__3165\ : InMux
    port map (
            O => \N__25495\,
            I => \ADC_IAC.n20678\
        );

    \I__3164\ : InMux
    port map (
            O => \N__25492\,
            I => \ADC_IAC.n20679\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__25489\,
            I => \N__25486\
        );

    \I__3162\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25483\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__25483\,
            I => n20_adj_1790
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__25480\,
            I => \n23498_cascade_\
        );

    \I__3159\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25473\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__25476\,
            I => \N__25470\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__25473\,
            I => \N__25467\
        );

    \I__3156\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25464\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__25467\,
            I => buf_adcdata_vdc_20
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__25464\,
            I => buf_adcdata_vdc_20
        );

    \I__3153\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25456\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25453\
        );

    \I__3151\ : Span4Mux_v
    port map (
            O => \N__25453\,
            I => \N__25450\
        );

    \I__3150\ : Sp12to4
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__3149\ : Span12Mux_h
    port map (
            O => \N__25447\,
            I => \N__25442\
        );

    \I__3148\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25439\
        );

    \I__3147\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25436\
        );

    \I__3146\ : Span12Mux_v
    port map (
            O => \N__25442\,
            I => \N__25433\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25428\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__25436\,
            I => \N__25428\
        );

    \I__3143\ : Odrv12
    port map (
            O => \N__25433\,
            I => buf_adcdata_vac_20
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__25428\,
            I => buf_adcdata_vac_20
        );

    \I__3141\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__25420\,
            I => n16_adj_1787
        );

    \I__3139\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__25414\,
            I => n17_adj_1788
        );

    \I__3137\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25408\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__25405\,
            I => n23540
        );

    \I__3134\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__3132\ : Span12Mux_s9_h
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__3131\ : Span12Mux_h
    port map (
            O => \N__25393\,
            I => \N__25389\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__25392\,
            I => \N__25385\
        );

    \I__3129\ : Span12Mux_v
    port map (
            O => \N__25389\,
            I => \N__25382\
        );

    \I__3128\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25377\
        );

    \I__3127\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25377\
        );

    \I__3126\ : Odrv12
    port map (
            O => \N__25382\,
            I => buf_adcdata_iac_23
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__25377\,
            I => buf_adcdata_iac_23
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__25372\,
            I => \N__25368\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__25371\,
            I => \N__25365\
        );

    \I__3122\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25360\
        );

    \I__3121\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25360\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__25360\,
            I => cmd_rdadctmp_31
        );

    \I__3119\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25351\
        );

    \I__3118\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25351\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__25351\,
            I => comm_test_buf_24_22
        );

    \I__3116\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25344\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__25347\,
            I => \N__25341\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25337\
        );

    \I__3113\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25334\
        );

    \I__3112\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25331\
        );

    \I__3111\ : Span4Mux_h
    port map (
            O => \N__25337\,
            I => \N__25328\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__25334\,
            I => buf_dds1_15
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__25331\,
            I => buf_dds1_15
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__25328\,
            I => buf_dds1_15
        );

    \I__3107\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25318\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__25318\,
            I => n111_adj_1771
        );

    \I__3105\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25312\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__25312\,
            I => \N__25308\
        );

    \I__3103\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25305\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__25308\,
            I => buf_adcdata_vdc_8
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__25305\,
            I => buf_adcdata_vdc_8
        );

    \I__3100\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__25297\,
            I => \N__25294\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__25294\,
            I => \N__25291\
        );

    \I__3097\ : Sp12to4
    port map (
            O => \N__25291\,
            I => \N__25287\
        );

    \I__3096\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25284\
        );

    \I__3095\ : Span12Mux_h
    port map (
            O => \N__25287\,
            I => \N__25280\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__25284\,
            I => \N__25277\
        );

    \I__3093\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25274\
        );

    \I__3092\ : Span12Mux_h
    port map (
            O => \N__25280\,
            I => \N__25271\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__25277\,
            I => \N__25268\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__25274\,
            I => buf_adcdata_vac_8
        );

    \I__3089\ : Odrv12
    port map (
            O => \N__25271\,
            I => buf_adcdata_vac_8
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__25268\,
            I => buf_adcdata_vac_8
        );

    \I__3087\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25258\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__25252\,
            I => n30_adj_1695
        );

    \I__3083\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25246\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__25243\,
            I => \N__25239\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__25242\,
            I => \N__25236\
        );

    \I__3079\ : Span4Mux_h
    port map (
            O => \N__25239\,
            I => \N__25233\
        );

    \I__3078\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25230\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__25233\,
            I => \buf_readRTD_11\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__25230\,
            I => \buf_readRTD_11\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__25225\,
            I => \N__25221\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__25224\,
            I => \N__25218\
        );

    \I__3073\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25212\
        );

    \I__3072\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25212\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__25217\,
            I => \N__25209\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25206\
        );

    \I__3069\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25203\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__25206\,
            I => \N__25198\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__25203\,
            I => \N__25198\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__25198\,
            I => \N__25193\
        );

    \I__3065\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25188\
        );

    \I__3064\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25188\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__25193\,
            I => \buf_cfgRTD_3\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__25188\,
            I => \buf_cfgRTD_3\
        );

    \I__3061\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25180\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25176\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__25179\,
            I => \N__25173\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__25176\,
            I => \N__25170\
        );

    \I__3057\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25167\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__25170\,
            I => buf_adcdata_vdc_6
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__25167\,
            I => buf_adcdata_vdc_6
        );

    \I__3054\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25159\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__25159\,
            I => \N__25155\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__25158\,
            I => \N__25152\
        );

    \I__3051\ : Span12Mux_s10_h
    port map (
            O => \N__25155\,
            I => \N__25149\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25146\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__25149\,
            I => buf_adcdata_vdc_22
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__25146\,
            I => buf_adcdata_vdc_22
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__3046\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25134\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \N__25131\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__25134\,
            I => \N__25128\
        );

    \I__3043\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25125\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__25128\,
            I => \N__25121\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__25125\,
            I => \N__25118\
        );

    \I__3040\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25115\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__25121\,
            I => cmd_rdadctmp_26_adj_1522
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__25118\,
            I => cmd_rdadctmp_26_adj_1522
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__25115\,
            I => cmd_rdadctmp_26_adj_1522
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__25108\,
            I => \n112_adj_1786_cascade_\
        );

    \I__3035\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25101\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__25104\,
            I => \N__25098\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__25101\,
            I => \N__25095\
        );

    \I__3032\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25092\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__25095\,
            I => buf_adcdata_vdc_10
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__25092\,
            I => buf_adcdata_vdc_10
        );

    \I__3029\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25084\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__25081\,
            I => \N__25078\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__25078\,
            I => \N__25073\
        );

    \I__3025\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25070\
        );

    \I__3024\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25067\
        );

    \I__3023\ : Sp12to4
    port map (
            O => \N__25073\,
            I => \N__25064\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__25070\,
            I => \N__25059\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25059\
        );

    \I__3020\ : Span12Mux_h
    port map (
            O => \N__25064\,
            I => \N__25056\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__25059\,
            I => buf_adcdata_vac_10
        );

    \I__3018\ : Odrv12
    port map (
            O => \N__25056\,
            I => buf_adcdata_vac_10
        );

    \I__3017\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25048\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__25048\,
            I => n19_adj_1747
        );

    \I__3015\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25041\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__25044\,
            I => \N__25038\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__25041\,
            I => \N__25035\
        );

    \I__3012\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25032\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__25035\,
            I => buf_adcdata_vdc_15
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__25032\,
            I => buf_adcdata_vdc_15
        );

    \I__3009\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25023\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__25026\,
            I => \N__25020\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__25023\,
            I => \N__25017\
        );

    \I__3006\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25014\
        );

    \I__3005\ : Odrv12
    port map (
            O => \N__25017\,
            I => buf_adcdata_vdc_7
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__25014\,
            I => buf_adcdata_vdc_7
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__3002\ : InMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24999\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__25002\,
            I => \N__24996\
        );

    \I__2999\ : Span12Mux_v
    port map (
            O => \N__24999\,
            I => \N__24993\
        );

    \I__2998\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24990\
        );

    \I__2997\ : Odrv12
    port map (
            O => \N__24993\,
            I => buf_adcdata_vdc_23
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__24990\,
            I => buf_adcdata_vdc_23
        );

    \I__2995\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24982\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__24982\,
            I => \N__24979\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__24979\,
            I => \N__24975\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__24978\,
            I => \N__24972\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__24975\,
            I => \N__24969\
        );

    \I__2990\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24966\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__24969\,
            I => buf_adcdata_vdc_4
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__24966\,
            I => buf_adcdata_vdc_4
        );

    \I__2987\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__24958\,
            I => \N__24954\
        );

    \I__2985\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24951\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__24954\,
            I => buf_adcdata_vdc_9
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__24951\,
            I => buf_adcdata_vdc_9
        );

    \I__2982\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__24943\,
            I => \RTD.n17\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__24940\,
            I => \N__24937\
        );

    \I__2979\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24930\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__24933\,
            I => \N__24925\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__24930\,
            I => \N__24919\
        );

    \I__2975\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24914\
        );

    \I__2974\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24914\
        );

    \I__2973\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24905\
        );

    \I__2972\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24905\
        );

    \I__2971\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24905\
        );

    \I__2970\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24905\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__24919\,
            I => \N__24902\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__24914\,
            I => \RTD.n79\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__24905\,
            I => \RTD.n79\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__24902\,
            I => \RTD.n79\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__2964\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__24889\,
            I => n12356
        );

    \I__2962\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N__24880\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__24880\,
            I => n22388
        );

    \I__2959\ : IoInMux
    port map (
            O => \N__24877\,
            I => \N__24874\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__2957\ : Span4Mux_s1_h
    port map (
            O => \N__24871\,
            I => \N__24868\
        );

    \I__2956\ : Span4Mux_h
    port map (
            O => \N__24868\,
            I => \N__24865\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__24865\,
            I => \N__24861\
        );

    \I__2954\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24858\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__24861\,
            I => \VDC_SCLK\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__24858\,
            I => \VDC_SCLK\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__24853\,
            I => \n21892_cascade_\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__24850\,
            I => \N__24847\
        );

    \I__2949\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24844\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__24844\,
            I => \N__24841\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__24841\,
            I => \N__24838\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__2945\ : IoSpan4Mux
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__24832\,
            I => \IAC_MISO\
        );

    \I__2943\ : IoInMux
    port map (
            O => \N__24829\,
            I => \N__24826\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24823\
        );

    \I__2941\ : Span12Mux_s6_v
    port map (
            O => \N__24823\,
            I => \N__24820\
        );

    \I__2940\ : Odrv12
    port map (
            O => \N__24820\,
            I => \GB_BUFFER_DDS_MCLK1_THRU_CO\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__2938\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24811\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__24811\,
            I => \CLK_DDS.tmp_buf_0\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24805\
        );

    \I__2935\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__24802\,
            I => \CLK_DDS.tmp_buf_1\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__24799\,
            I => \N__24796\
        );

    \I__2932\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24793\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__24793\,
            I => \CLK_DDS.tmp_buf_2\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__2929\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24784\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__24784\,
            I => \CLK_DDS.tmp_buf_3\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__24781\,
            I => \N__24778\
        );

    \I__2926\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24775\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__24775\,
            I => \CLK_DDS.tmp_buf_4\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__2923\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__24766\,
            I => \CLK_DDS.tmp_buf_5\
        );

    \I__2921\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24731\
        );

    \I__2920\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24731\
        );

    \I__2919\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24731\
        );

    \I__2918\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24731\
        );

    \I__2917\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24731\
        );

    \I__2916\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24731\
        );

    \I__2915\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24731\
        );

    \I__2914\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24731\
        );

    \I__2913\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24714\
        );

    \I__2912\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24714\
        );

    \I__2911\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24714\
        );

    \I__2910\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24714\
        );

    \I__2909\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24714\
        );

    \I__2908\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24714\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24714\
        );

    \I__2906\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24714\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24711\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24708\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__24711\,
            I => \N__24698\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__24708\,
            I => \N__24698\
        );

    \I__2901\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24695\
        );

    \I__2900\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24692\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__24705\,
            I => \N__24685\
        );

    \I__2898\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24679\
        );

    \I__2897\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24679\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__24698\,
            I => \N__24672\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__24695\,
            I => \N__24672\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__24692\,
            I => \N__24672\
        );

    \I__2893\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24669\
        );

    \I__2892\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24666\
        );

    \I__2891\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24663\
        );

    \I__2890\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24656\
        );

    \I__2889\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24656\
        );

    \I__2888\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24656\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__24679\,
            I => \N__24647\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__24672\,
            I => \N__24647\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24647\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__24666\,
            I => \N__24647\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__24663\,
            I => dds_state_2_adj_1508
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__24656\,
            I => dds_state_2_adj_1508
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__24647\,
            I => dds_state_2_adj_1508
        );

    \I__2880\ : CEMux
    port map (
            O => \N__24640\,
            I => \N__24636\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__24639\,
            I => \N__24615\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__24636\,
            I => \N__24606\
        );

    \I__2877\ : SRMux
    port map (
            O => \N__24635\,
            I => \N__24603\
        );

    \I__2876\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24588\
        );

    \I__2875\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24588\
        );

    \I__2874\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24588\
        );

    \I__2873\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24588\
        );

    \I__2872\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24588\
        );

    \I__2871\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24588\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24588\
        );

    \I__2869\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24585\
        );

    \I__2868\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24568\
        );

    \I__2867\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24568\
        );

    \I__2866\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24568\
        );

    \I__2865\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24568\
        );

    \I__2864\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24568\
        );

    \I__2863\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24568\
        );

    \I__2862\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24568\
        );

    \I__2861\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24568\
        );

    \I__2860\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24565\
        );

    \I__2859\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24560\
        );

    \I__2858\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24560\
        );

    \I__2857\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24557\
        );

    \I__2856\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24550\
        );

    \I__2855\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24550\
        );

    \I__2854\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24550\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__24609\,
            I => \N__24547\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__24606\,
            I => \N__24543\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24540\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24537\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24530\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24530\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24530\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__24560\,
            I => \N__24523\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__24557\,
            I => \N__24523\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24523\
        );

    \I__2843\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24519\
        );

    \I__2842\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24516\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__24543\,
            I => \N__24507\
        );

    \I__2840\ : Span4Mux_v
    port map (
            O => \N__24540\,
            I => \N__24507\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__24537\,
            I => \N__24507\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__24530\,
            I => \N__24507\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__24523\,
            I => \N__24504\
        );

    \I__2836\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24501\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__24519\,
            I => \N__24496\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24496\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__24507\,
            I => dds_state_1_adj_1509
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__24504\,
            I => dds_state_1_adj_1509
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__24501\,
            I => dds_state_1_adj_1509
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__24496\,
            I => dds_state_1_adj_1509
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__2828\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__24481\,
            I => \CLK_DDS.tmp_buf_6\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__2825\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24472\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__24472\,
            I => \CLK_DDS.tmp_buf_7\
        );

    \I__2823\ : CEMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24462\
        );

    \I__2821\ : CEMux
    port map (
            O => \N__24465\,
            I => \N__24459\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__24462\,
            I => \N__24456\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24453\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__24456\,
            I => \N__24450\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__24453\,
            I => \N__24447\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__24450\,
            I => \N__24442\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__24447\,
            I => \N__24442\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__24439\,
            I => \CLK_DDS.n13376\
        );

    \I__2812\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24433\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__24433\,
            I => n19_adj_1765
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__2809\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24424\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__2807\ : Span12Mux_v
    port map (
            O => \N__24421\,
            I => \N__24418\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__24418\,
            I => n20_adj_1766
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__24415\,
            I => \N__24412\
        );

    \I__2804\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__24409\,
            I => \CLK_DDS.tmp_buf_10\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__24406\,
            I => \N__24403\
        );

    \I__2801\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__24400\,
            I => \CLK_DDS.tmp_buf_11\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__24397\,
            I => \N__24394\
        );

    \I__2798\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__24391\,
            I => \CLK_DDS.tmp_buf_12\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__2795\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__24382\,
            I => \CLK_DDS.tmp_buf_13\
        );

    \I__2793\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__24376\,
            I => \CLK_DDS.tmp_buf_14\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__2790\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24367\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__24367\,
            I => \CLK_DDS.tmp_buf_9\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__2787\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__24358\,
            I => \CLK_DDS.tmp_buf_8\
        );

    \I__2785\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24351\
        );

    \I__2784\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24348\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__24351\,
            I => tmp_buf_15_adj_1511
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__24348\,
            I => tmp_buf_15_adj_1511
        );

    \I__2781\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24336\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__24339\,
            I => \N__24333\
        );

    \I__2778\ : Span4Mux_v
    port map (
            O => \N__24336\,
            I => \N__24330\
        );

    \I__2777\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24327\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__24330\,
            I => \buf_readRTD_2\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__24327\,
            I => \buf_readRTD_2\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__24322\,
            I => \N__24318\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__24321\,
            I => \N__24315\
        );

    \I__2772\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24312\
        );

    \I__2771\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24309\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__24312\,
            I => \N__24306\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__24309\,
            I => \N__24302\
        );

    \I__2768\ : Span12Mux_s9_h
    port map (
            O => \N__24306\,
            I => \N__24299\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24296\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__24302\,
            I => cmd_rdadctmp_12_adj_1536
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__24299\,
            I => cmd_rdadctmp_12_adj_1536
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__24296\,
            I => cmd_rdadctmp_12_adj_1536
        );

    \I__2763\ : IoInMux
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__2761\ : Span4Mux_s3_v
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__24280\,
            I => \N__24277\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__24274\,
            I => \N__24270\
        );

    \I__2757\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24267\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__24270\,
            I => \DDS_MOSI1\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__24267\,
            I => \DDS_MOSI1\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__2753\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24255\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__24258\,
            I => \N__24252\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24249\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24245\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__24249\,
            I => \N__24242\
        );

    \I__2748\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24239\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24245\,
            I => cmd_rdadctmp_22_adj_1526
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__24242\,
            I => cmd_rdadctmp_22_adj_1526
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__24239\,
            I => cmd_rdadctmp_22_adj_1526
        );

    \I__2744\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24229\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24225\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__24228\,
            I => \N__24222\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__24225\,
            I => \N__24219\
        );

    \I__2740\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24215\
        );

    \I__2739\ : Sp12to4
    port map (
            O => \N__24219\,
            I => \N__24212\
        );

    \I__2738\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24209\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24204\
        );

    \I__2736\ : Span12Mux_h
    port map (
            O => \N__24212\,
            I => \N__24204\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__24209\,
            I => buf_adcdata_vac_15
        );

    \I__2734\ : Odrv12
    port map (
            O => \N__24204\,
            I => buf_adcdata_vac_15
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \n19_adj_1714_cascade_\
        );

    \I__2732\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24193\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N__24189\
        );

    \I__2730\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24186\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__24189\,
            I => \buf_readRTD_7\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__24186\,
            I => \buf_readRTD_7\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__24181\,
            I => \N__24177\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24172\
        );

    \I__2725\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24172\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__24172\,
            I => \RTD.adress_2\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__24169\,
            I => \N__24166\
        );

    \I__2722\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24163\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__24163\,
            I => \RTD.adress_0\
        );

    \I__2720\ : CEMux
    port map (
            O => \N__24160\,
            I => \N__24151\
        );

    \I__2719\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24138\
        );

    \I__2718\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24138\
        );

    \I__2717\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24138\
        );

    \I__2716\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24138\
        );

    \I__2715\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24138\
        );

    \I__2714\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24138\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__24151\,
            I => \RTD.n13441\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__24138\,
            I => \RTD.n13441\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__24133\,
            I => \N__24129\
        );

    \I__2710\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24126\
        );

    \I__2709\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24123\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__24126\,
            I => \RTD.adress_1\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__24123\,
            I => \RTD.adress_1\
        );

    \I__2706\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24115\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24111\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__24114\,
            I => \N__24108\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__24111\,
            I => \N__24104\
        );

    \I__2702\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24101\
        );

    \I__2701\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24098\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__24104\,
            I => read_buf_6
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__24101\,
            I => read_buf_6
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__24098\,
            I => read_buf_6
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__24091\,
            I => \N__24084\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__24090\,
            I => \N__24080\
        );

    \I__2695\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24073\
        );

    \I__2694\ : InMux
    port map (
            O => \N__24088\,
            I => \N__24068\
        );

    \I__2693\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24068\
        );

    \I__2692\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24062\
        );

    \I__2691\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24062\
        );

    \I__2690\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24055\
        );

    \I__2689\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24055\
        );

    \I__2688\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24055\
        );

    \I__2687\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24049\
        );

    \I__2686\ : InMux
    port map (
            O => \N__24076\,
            I => \N__24046\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__24073\,
            I => \N__24041\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24041\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__24067\,
            I => \N__24038\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__24062\,
            I => \N__24032\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__24055\,
            I => \N__24032\
        );

    \I__2680\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24027\
        );

    \I__2679\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24027\
        );

    \I__2678\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24024\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24019\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__24046\,
            I => \N__24019\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__24041\,
            I => \N__24016\
        );

    \I__2674\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24013\
        );

    \I__2673\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24010\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__24032\,
            I => \N__24007\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__24027\,
            I => \N__24004\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__23999\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__24019\,
            I => \N__23999\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__24016\,
            I => n21989
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__24013\,
            I => n21989
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__24010\,
            I => n21989
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__24007\,
            I => n21989
        );

    \I__2664\ : Odrv12
    port map (
            O => \N__24004\,
            I => n21989
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__23999\,
            I => n21989
        );

    \I__2662\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23967\
        );

    \I__2661\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23967\
        );

    \I__2660\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23967\
        );

    \I__2659\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23960\
        );

    \I__2658\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23960\
        );

    \I__2657\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23960\
        );

    \I__2656\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23955\
        );

    \I__2655\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23955\
        );

    \I__2654\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23950\
        );

    \I__2653\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23950\
        );

    \I__2652\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23945\
        );

    \I__2651\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23945\
        );

    \I__2650\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23942\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__23967\,
            I => \N__23934\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23934\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__23955\,
            I => \N__23931\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__23950\,
            I => \N__23928\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23925\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23922\
        );

    \I__2643\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23915\
        );

    \I__2642\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23915\
        );

    \I__2641\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23915\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__23934\,
            I => \N__23912\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__23931\,
            I => \N__23907\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__23928\,
            I => \N__23907\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__23925\,
            I => \N__23902\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__23922\,
            I => \N__23902\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__23915\,
            I => n13584
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__23912\,
            I => n13584
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__23907\,
            I => n13584
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__23902\,
            I => n13584
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23888\
        );

    \I__2630\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23881\
        );

    \I__2629\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23881\
        );

    \I__2628\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23881\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__23881\,
            I => read_buf_7
        );

    \I__2626\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__23875\,
            I => \N__23872\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__23872\,
            I => \N__23869\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__23869\,
            I => \N__23865\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__23868\,
            I => \N__23862\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__23865\,
            I => \N__23858\
        );

    \I__2620\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23855\
        );

    \I__2619\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23852\
        );

    \I__2618\ : Sp12to4
    port map (
            O => \N__23858\,
            I => \N__23849\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__23855\,
            I => buf_adcdata_vac_9
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__23852\,
            I => buf_adcdata_vac_9
        );

    \I__2615\ : Odrv12
    port map (
            O => \N__23849\,
            I => buf_adcdata_vac_9
        );

    \I__2614\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__23839\,
            I => n19_adj_1752
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23831\
        );

    \I__2611\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23828\
        );

    \I__2610\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23823\
        );

    \I__2609\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23823\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__23828\,
            I => read_buf_8
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__23823\,
            I => read_buf_8
        );

    \I__2606\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23807\
        );

    \I__2605\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23804\
        );

    \I__2604\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23799\
        );

    \I__2603\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23799\
        );

    \I__2602\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23796\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \N__23793\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__23812\,
            I => \N__23789\
        );

    \I__2599\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23784\
        );

    \I__2598\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23784\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23772\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23772\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__23799\,
            I => \N__23772\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__23796\,
            I => \N__23769\
        );

    \I__2593\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23764\
        );

    \I__2592\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23764\
        );

    \I__2591\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23761\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23758\
        );

    \I__2589\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23749\
        );

    \I__2588\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23749\
        );

    \I__2587\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23749\
        );

    \I__2586\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23749\
        );

    \I__2585\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23746\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__23772\,
            I => \N__23741\
        );

    \I__2583\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23741\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__23764\,
            I => \N__23736\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__23761\,
            I => \N__23736\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__23758\,
            I => \N__23733\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__23749\,
            I => n13603
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__23746\,
            I => n13603
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__23741\,
            I => n13603
        );

    \I__2576\ : Odrv12
    port map (
            O => \N__23736\,
            I => n13603
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__23733\,
            I => n13603
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__23722\,
            I => \N__23719\
        );

    \I__2573\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23711\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__23715\,
            I => \N__23708\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__23714\,
            I => \N__23705\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__23711\,
            I => \N__23702\
        );

    \I__2568\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23699\
        );

    \I__2567\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23696\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__23702\,
            I => read_buf_9
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__23699\,
            I => read_buf_9
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__23696\,
            I => read_buf_9
        );

    \I__2563\ : InMux
    port map (
            O => \N__23689\,
            I => \N__23682\
        );

    \I__2562\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23679\
        );

    \I__2561\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23675\
        );

    \I__2560\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23670\
        );

    \I__2559\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23670\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23667\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23664\
        );

    \I__2556\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23661\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__23675\,
            I => \RTD.adress_7_N_1009_7\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__23670\,
            I => \RTD.adress_7_N_1009_7\
        );

    \I__2553\ : Odrv12
    port map (
            O => \N__23667\,
            I => \RTD.adress_7_N_1009_7\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__23664\,
            I => \RTD.adress_7_N_1009_7\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__23661\,
            I => \RTD.adress_7_N_1009_7\
        );

    \I__2550\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23645\
        );

    \I__2549\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23640\
        );

    \I__2548\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23640\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__23645\,
            I => \RTD.n11\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__23640\,
            I => \RTD.n11\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__23635\,
            I => \RTD.n11_cascade_\
        );

    \I__2544\ : CEMux
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__23623\,
            I => \RTD.n13488\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__23620\,
            I => \RTD.n13488_cascade_\
        );

    \I__2539\ : SRMux
    port map (
            O => \N__23617\,
            I => \N__23614\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__23608\,
            I => \RTD.n15585\
        );

    \I__2535\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23602\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__23602\,
            I => \RTD.n22081\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__23599\,
            I => \N__23595\
        );

    \I__2532\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23592\
        );

    \I__2531\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__23592\,
            I => \RTD.adress_6\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__23589\,
            I => \RTD.adress_6\
        );

    \I__2528\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23578\
        );

    \I__2527\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23578\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__23578\,
            I => \RTD.adress_5\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__23575\,
            I => \N__23571\
        );

    \I__2524\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23566\
        );

    \I__2523\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23566\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__23566\,
            I => \RTD.adress_4\
        );

    \I__2521\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23557\
        );

    \I__2520\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23557\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__23557\,
            I => \RTD.adress_3\
        );

    \I__2518\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__2517\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23548\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__23548\,
            I => \RTD.cfg_buf_6\
        );

    \I__2515\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23539\
        );

    \I__2514\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23539\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__23539\,
            I => \RTD.cfg_buf_5\
        );

    \I__2512\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__23533\,
            I => \RTD.n12\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__2509\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23523\
        );

    \I__2508\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23520\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__23523\,
            I => \RTD.cfg_buf_1\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__23520\,
            I => \RTD.cfg_buf_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23512\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__23512\,
            I => \RTD.n20093\
        );

    \I__2503\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23499\
        );

    \I__2502\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23492\
        );

    \I__2501\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23492\
        );

    \I__2500\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23492\
        );

    \I__2499\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23483\
        );

    \I__2498\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23483\
        );

    \I__2497\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23483\
        );

    \I__2496\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23483\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__23499\,
            I => \RTD.n13482\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__23492\,
            I => \RTD.n13482\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__23483\,
            I => \RTD.n13482\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__23476\,
            I => \N__23471\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__23475\,
            I => \N__23468\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__23474\,
            I => \N__23465\
        );

    \I__2489\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23455\
        );

    \I__2488\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23446\
        );

    \I__2487\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23446\
        );

    \I__2486\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23446\
        );

    \I__2485\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23446\
        );

    \I__2484\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23443\
        );

    \I__2483\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23436\
        );

    \I__2482\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23436\
        );

    \I__2481\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23436\
        );

    \I__2480\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23433\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23428\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__23446\,
            I => \N__23428\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__23443\,
            I => \N__23425\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__23436\,
            I => \RTD.n68\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__23433\,
            I => \RTD.n68\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__23428\,
            I => \RTD.n68\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__23425\,
            I => \RTD.n68\
        );

    \I__2472\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23412\
        );

    \I__2471\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23409\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__23412\,
            I => \RTD.cfg_buf_7\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__23409\,
            I => \RTD.cfg_buf_7\
        );

    \I__2468\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23400\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__23403\,
            I => \N__23397\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__23400\,
            I => \N__23394\
        );

    \I__2465\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23391\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__23394\,
            I => \buf_readRTD_14\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__23391\,
            I => \buf_readRTD_14\
        );

    \I__2462\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23380\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__23380\,
            I => \RTD.n68_adj_1498\
        );

    \I__2459\ : CEMux
    port map (
            O => \N__23377\,
            I => \N__23374\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__23371\,
            I => \N__23368\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__23368\,
            I => \RTD.n21954\
        );

    \I__2455\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23360\
        );

    \I__2454\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23357\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \N__23354\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23349\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__23357\,
            I => \N__23349\
        );

    \I__2450\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23346\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__23349\,
            I => \N__23342\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23339\
        );

    \I__2447\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23336\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__23342\,
            I => \N__23333\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__23339\,
            I => \N__23328\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23328\
        );

    \I__2443\ : Span4Mux_h
    port map (
            O => \N__23333\,
            I => \N__23325\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__23328\,
            I => \N__23322\
        );

    \I__2441\ : Sp12to4
    port map (
            O => \N__23325\,
            I => \N__23317\
        );

    \I__2440\ : Sp12to4
    port map (
            O => \N__23322\,
            I => \N__23317\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__23317\,
            I => \RTD_DRDY\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__23314\,
            I => \RTD.n21954_cascade_\
        );

    \I__2437\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23308\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__23308\,
            I => \RTD.n21955\
        );

    \I__2435\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23302\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__23302\,
            I => \RTD.n21988\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__23299\,
            I => \RTD.n7_adj_1497_cascade_\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__23296\,
            I => \n13603_cascade_\
        );

    \I__2431\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23288\
        );

    \I__2430\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23283\
        );

    \I__2429\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23283\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__23288\,
            I => read_buf_5
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__23283\,
            I => read_buf_5
        );

    \I__2426\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23275\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__23275\,
            I => \RTD.n62\
        );

    \I__2424\ : CEMux
    port map (
            O => \N__23272\,
            I => \N__23268\
        );

    \I__2423\ : CEMux
    port map (
            O => \N__23271\,
            I => \N__23265\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__23268\,
            I => \RTD.n12274\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__23265\,
            I => \RTD.n12274\
        );

    \I__2420\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23257\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__23257\,
            I => \RTD.n11_adj_1500\
        );

    \I__2418\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23251\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23247\
        );

    \I__2416\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23244\
        );

    \I__2415\ : Span12Mux_s11_h
    port map (
            O => \N__23247\,
            I => \N__23241\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__23244\,
            I => \N__23238\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__23241\,
            I => \N__23234\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__23238\,
            I => \N__23231\
        );

    \I__2411\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23228\
        );

    \I__2410\ : Span12Mux_h
    port map (
            O => \N__23234\,
            I => \N__23225\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__23231\,
            I => \N__23222\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__23228\,
            I => buf_adcdata_vac_23
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__23225\,
            I => buf_adcdata_vac_23
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__23222\,
            I => buf_adcdata_vac_23
        );

    \I__2405\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__2403\ : Span12Mux_v
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__2402\ : Odrv12
    port map (
            O => \N__23206\,
            I => n23435
        );

    \I__2401\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23197\
        );

    \I__2400\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23194\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23191\
        );

    \I__2398\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23188\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__23197\,
            I => \N__23185\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23182\
        );

    \I__2395\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23179\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23176\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__23185\,
            I => \N__23173\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__23182\,
            I => \N__23170\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__23179\,
            I => \RTD.mode\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__23176\,
            I => \RTD.mode\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__23173\,
            I => \RTD.mode\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__23170\,
            I => \RTD.mode\
        );

    \I__2387\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23155\
        );

    \I__2386\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23155\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__23155\,
            I => cmd_rdadctmp_31_adj_1517
        );

    \I__2384\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__23149\,
            I => \N__23146\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__23146\,
            I => \N__23142\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__23145\,
            I => \N__23139\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__23142\,
            I => \N__23135\
        );

    \I__2379\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23130\
        );

    \I__2378\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23130\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__23135\,
            I => cmd_rdadctmp_29_adj_1519
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__23130\,
            I => cmd_rdadctmp_29_adj_1519
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__23125\,
            I => \N__23120\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__23124\,
            I => \N__23117\
        );

    \I__2373\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23110\
        );

    \I__2372\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23110\
        );

    \I__2371\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23110\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__23110\,
            I => cmd_rdadctmp_30_adj_1518
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__23107\,
            I => \n21948_cascade_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__2365\ : Sp12to4
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__2364\ : Span12Mux_v
    port map (
            O => \N__23092\,
            I => \N__23088\
        );

    \I__2363\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23084\
        );

    \I__2362\ : Span12Mux_h
    port map (
            O => \N__23088\,
            I => \N__23081\
        );

    \I__2361\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23078\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__23084\,
            I => buf_adcdata_vac_22
        );

    \I__2359\ : Odrv12
    port map (
            O => \N__23081\,
            I => buf_adcdata_vac_22
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__23078\,
            I => buf_adcdata_vac_22
        );

    \I__2357\ : IoInMux
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23065\
        );

    \I__2355\ : IoSpan4Mux
    port map (
            O => \N__23065\,
            I => \N__23062\
        );

    \I__2354\ : Span4Mux_s3_v
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__23059\,
            I => \N__23056\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__23056\,
            I => \AC_ADC_SYNC\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__23053\,
            I => \N__23049\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23044\
        );

    \I__2349\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23044\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23041\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__23041\,
            I => \N__23037\
        );

    \I__2346\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23034\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__23037\,
            I => cmd_rdadctmp_23_adj_1525
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__23034\,
            I => cmd_rdadctmp_23_adj_1525
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__2342\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__23023\,
            I => \N__23018\
        );

    \I__2340\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23013\
        );

    \I__2339\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23013\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__23018\,
            I => cmd_rdadctmp_24_adj_1524
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__23013\,
            I => cmd_rdadctmp_24_adj_1524
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__2335\ : InMux
    port map (
            O => \N__23005\,
            I => \N__23001\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \N__22998\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22995\
        );

    \I__2332\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22991\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__22995\,
            I => \N__22988\
        );

    \I__2330\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22985\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__22991\,
            I => cmd_rdadctmp_28_adj_1520
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__22988\,
            I => cmd_rdadctmp_28_adj_1520
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__22985\,
            I => cmd_rdadctmp_28_adj_1520
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__2325\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__22972\,
            I => \N__22969\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__22969\,
            I => \N__22964\
        );

    \I__2322\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22959\
        );

    \I__2321\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22959\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__22964\,
            I => cmd_rdadctmp_15
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__22959\,
            I => cmd_rdadctmp_15
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__2317\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22947\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__22950\,
            I => \N__22944\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22940\
        );

    \I__2314\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22935\
        );

    \I__2313\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22935\
        );

    \I__2312\ : Odrv12
    port map (
            O => \N__22940\,
            I => cmd_rdadctmp_13_adj_1535
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__22935\,
            I => cmd_rdadctmp_13_adj_1535
        );

    \I__2310\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22922\
        );

    \I__2308\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22919\
        );

    \I__2307\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22916\
        );

    \I__2306\ : Span12Mux_v
    port map (
            O => \N__22922\,
            I => \N__22913\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__22919\,
            I => \N__22910\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__22916\,
            I => buf_adcdata_vac_5
        );

    \I__2303\ : Odrv12
    port map (
            O => \N__22913\,
            I => buf_adcdata_vac_5
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__22910\,
            I => buf_adcdata_vac_5
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__22903\,
            I => \N__22900\
        );

    \I__2300\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22892\
        );

    \I__2298\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22887\
        );

    \I__2297\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22887\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__22892\,
            I => cmd_rdadctmp_17_adj_1531
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__22887\,
            I => cmd_rdadctmp_17_adj_1531
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__22882\,
            I => \N__22878\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__22881\,
            I => \N__22875\
        );

    \I__2292\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22870\
        );

    \I__2291\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22870\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__22870\,
            I => \N__22866\
        );

    \I__2289\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__2288\ : Odrv12
    port map (
            O => \N__22866\,
            I => cmd_rdadctmp_18_adj_1530
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__22863\,
            I => cmd_rdadctmp_18_adj_1530
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__22858\,
            I => \n23543_cascade_\
        );

    \I__2285\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22849\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__22849\,
            I => n19_adj_1696
        );

    \I__2282\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22840\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__22837\,
            I => buf_data_iac_7
        );

    \I__2278\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__22825\,
            I => n22_adj_1691
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__2273\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22815\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__22818\,
            I => \N__22812\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22809\
        );

    \I__2270\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22805\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__22809\,
            I => \N__22802\
        );

    \I__2268\ : InMux
    port map (
            O => \N__22808\,
            I => \N__22799\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__22805\,
            I => cmd_rdadctmp_16_adj_1532
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__22802\,
            I => cmd_rdadctmp_16_adj_1532
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__22799\,
            I => cmd_rdadctmp_16_adj_1532
        );

    \I__2264\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__22789\,
            I => \RTD.cfg_tmp_3\
        );

    \I__2262\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__22783\,
            I => \RTD.cfg_tmp_4\
        );

    \I__2260\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__22777\,
            I => \RTD.cfg_tmp_5\
        );

    \I__2258\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__22771\,
            I => \RTD.cfg_tmp_6\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__2255\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__2253\ : Span4Mux_v
    port map (
            O => \N__22759\,
            I => \N__22755\
        );

    \I__2252\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22752\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__22755\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__22752\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2249\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__22744\,
            I => \N__22741\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__22741\,
            I => \N__22738\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__22738\,
            I => buf_data_iac_6
        );

    \I__2245\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22729\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__22729\,
            I => n22_adj_1694
        );

    \I__2242\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22719\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__22722\,
            I => \N__22716\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__22719\,
            I => \N__22713\
        );

    \I__2238\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22710\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__22713\,
            I => \buf_readRTD_1\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__22710\,
            I => \buf_readRTD_1\
        );

    \I__2235\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22702\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__22699\,
            I => \N__22695\
        );

    \I__2232\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22692\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__22695\,
            I => cmd_rdadctmp_2_adj_1546
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__22692\,
            I => cmd_rdadctmp_2_adj_1546
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__22687\,
            I => \N__22683\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__22686\,
            I => \N__22680\
        );

    \I__2227\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__2226\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22674\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__22677\,
            I => \N__22671\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22665\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__2222\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22662\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__22665\,
            I => cmd_rdadctmp_12
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__22662\,
            I => cmd_rdadctmp_12
        );

    \I__2219\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22650\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__22653\,
            I => \N__22647\
        );

    \I__2216\ : Span4Mux_v
    port map (
            O => \N__22650\,
            I => \N__22644\
        );

    \I__2215\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22641\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__22644\,
            I => \N__22638\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__22641\,
            I => \RTD.adress_7\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__22638\,
            I => \RTD.adress_7\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \RTD.n19_cascade_\
        );

    \I__2210\ : SRMux
    port map (
            O => \N__22630\,
            I => \N__22627\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__22627\,
            I => \RTD.n15396\
        );

    \I__2208\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22621\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__22621\,
            I => \RTD.n1\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__22618\,
            I => \RTD.n1_cascade_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22612\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__22612\,
            I => \RTD.cfg_tmp_0\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__22609\,
            I => \N__22606\
        );

    \I__2202\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22603\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__22603\,
            I => \RTD.cfg_tmp_1\
        );

    \I__2200\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__22597\,
            I => \RTD.cfg_tmp_2\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__22594\,
            I => \RTD.n68_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22585\
        );

    \I__2196\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22585\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__22585\,
            I => \RTD.cfg_buf_4\
        );

    \I__2194\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22576\
        );

    \I__2193\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22576\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__22576\,
            I => \RTD.cfg_buf_2\
        );

    \I__2191\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22567\
        );

    \I__2190\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22567\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__22567\,
            I => \RTD.cfg_buf_0\
        );

    \I__2188\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22561\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__22561\,
            I => \RTD.n10\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__22558\,
            I => \RTD.n9_cascade_\
        );

    \I__2185\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22549\
        );

    \I__2184\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22549\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__22549\,
            I => \RTD.cfg_buf_3\
        );

    \I__2182\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22540\
        );

    \I__2181\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22540\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__22540\,
            I => \RTD.n20051\
        );

    \I__2179\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__22531\,
            I => \N__22526\
        );

    \I__2176\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22521\
        );

    \I__2175\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22521\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__22526\,
            I => read_buf_0
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__22521\,
            I => read_buf_0
        );

    \I__2172\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22512\
        );

    \I__2171\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22509\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__22512\,
            I => \N__22503\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__22509\,
            I => \N__22503\
        );

    \I__2168\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22500\
        );

    \I__2167\ : Odrv12
    port map (
            O => \N__22503\,
            I => \RTD.read_buf_4\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__22500\,
            I => \RTD.read_buf_4\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__22495\,
            I => \n21989_cascade_\
        );

    \I__2164\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22486\
        );

    \I__2163\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22486\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22483\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__22483\,
            I => \N__22479\
        );

    \I__2160\ : InMux
    port map (
            O => \N__22482\,
            I => \N__22476\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__22479\,
            I => read_buf_1
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__22476\,
            I => read_buf_1
        );

    \I__2157\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__22468\,
            I => \N__22464\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__22467\,
            I => \N__22460\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__22464\,
            I => \N__22457\
        );

    \I__2153\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22452\
        );

    \I__2152\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22452\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__22457\,
            I => read_buf_2
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__22452\,
            I => read_buf_2
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__22447\,
            I => \RTD.n20051_cascade_\
        );

    \I__2148\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22441\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__22435\,
            I => \RTD.n22079\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__22432\,
            I => \RTD.n22599_cascade_\
        );

    \I__2143\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22425\
        );

    \I__2142\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22422\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__22425\,
            I => \N__22419\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__22422\,
            I => \RTD.n23689\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__22419\,
            I => \RTD.n23689\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__22414\,
            I => \RTD.n56_cascade_\
        );

    \I__2137\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__22405\,
            I => \RTD.n5\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__22399\,
            I => \RTD.n71\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__22396\,
            I => \RTD.n71_cascade_\
        );

    \I__2131\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__22390\,
            I => \RTD.n22623\
        );

    \I__2129\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22383\
        );

    \I__2128\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22380\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__22383\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__22380\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__2125\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22371\
        );

    \I__2124\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22368\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__22371\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__22368\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \ADC_VAC.n22109_cascade_\
        );

    \I__2120\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22356\
        );

    \I__2119\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22353\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__22356\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__22353\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__22348\,
            I => \ADC_VAC.n22126_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22341\
        );

    \I__2114\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22338\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__22341\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__22338\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__22333\,
            I => \ADC_VAC.n22389_cascade_\
        );

    \I__2110\ : CEMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__22324\,
            I => \ADC_VAC.n22030\
        );

    \I__2107\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__22318\,
            I => \ADC_VAC.n17\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__22315\,
            I => \N__22312\
        );

    \I__2104\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22307\
        );

    \I__2103\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22304\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22301\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22296\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__22304\,
            I => \N__22296\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__22301\,
            I => \N__22291\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__22296\,
            I => \N__22288\
        );

    \I__2097\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22283\
        );

    \I__2096\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22283\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__22291\,
            I => \N__22280\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__22288\,
            I => \N__22275\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__22283\,
            I => \N__22275\
        );

    \I__2092\ : Span4Mux_h
    port map (
            O => \N__22280\,
            I => \N__22272\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__22275\,
            I => \VAC_DRDY\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__22272\,
            I => \VAC_DRDY\
        );

    \I__2089\ : CEMux
    port map (
            O => \N__22267\,
            I => \N__22263\
        );

    \I__2088\ : CEMux
    port map (
            O => \N__22266\,
            I => \N__22260\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22257\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__22260\,
            I => \N__22254\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__22257\,
            I => \N__22251\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__22254\,
            I => \N__22248\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__22251\,
            I => \ADC_VAC.n12\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__22248\,
            I => \ADC_VAC.n12\
        );

    \I__2081\ : IoInMux
    port map (
            O => \N__22243\,
            I => \N__22240\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__2079\ : Span12Mux_s8_h
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__22234\,
            I => \RTD_CS\
        );

    \I__2077\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__22228\,
            I => \RTD.n22382\
        );

    \I__2075\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__22222\,
            I => n22_adj_1697
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__22219\,
            I => \N__22216\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22213\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__22213\,
            I => \N__22209\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__22212\,
            I => \N__22206\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__22209\,
            I => \N__22202\
        );

    \I__2068\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22199\
        );

    \I__2067\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22196\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__22202\,
            I => cmd_rdadctmp_15_adj_1533
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__22199\,
            I => cmd_rdadctmp_15_adj_1533
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__22196\,
            I => cmd_rdadctmp_15_adj_1533
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__2062\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22182\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__22185\,
            I => \N__22179\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__22182\,
            I => \N__22175\
        );

    \I__2059\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22170\
        );

    \I__2058\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22170\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__22175\,
            I => cmd_rdadctmp_13
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__22170\,
            I => cmd_rdadctmp_13
        );

    \I__2055\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__22162\,
            I => \N__22158\
        );

    \I__2053\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22154\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__22158\,
            I => \N__22151\
        );

    \I__2051\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22148\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__22154\,
            I => buf_adcdata_iac_5
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__22151\,
            I => buf_adcdata_iac_5
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__22148\,
            I => buf_adcdata_iac_5
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__22141\,
            I => \ADC_VAC.n13747_cascade_\
        );

    \I__2046\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__22135\,
            I => \ADC_VAC.n13842\
        );

    \I__2044\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22128\
        );

    \I__2043\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22125\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__22128\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__22125\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__2040\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22116\
        );

    \I__2039\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22113\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__22116\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__22113\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__22108\,
            I => \N__22104\
        );

    \I__2035\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22101\
        );

    \I__2034\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22098\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__22101\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__22098\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__2031\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22089\
        );

    \I__2030\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22086\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__22089\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__22086\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__2027\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22075\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__22072\,
            I => buf_data_iac_5
        );

    \I__2023\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__22066\,
            I => \N__22063\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__22063\,
            I => \N__22058\
        );

    \I__2020\ : InMux
    port map (
            O => \N__22062\,
            I => \N__22053\
        );

    \I__2019\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22053\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__22058\,
            I => buf_adcdata_iac_6
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__22053\,
            I => buf_adcdata_iac_6
        );

    \I__2016\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__22045\,
            I => \N__22041\
        );

    \I__2014\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22037\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__22041\,
            I => \N__22034\
        );

    \I__2012\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22031\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__22037\,
            I => buf_adcdata_iac_7
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__22034\,
            I => buf_adcdata_iac_7
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__22031\,
            I => buf_adcdata_iac_7
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__2007\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22012\
        );

    \I__2006\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22012\
        );

    \I__2005\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22012\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__22012\,
            I => cmd_rdadctmp_14
        );

    \I__2003\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__22006\,
            I => n19_adj_1700
        );

    \I__2001\ : InMux
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__21994\,
            I => buf_data_iac_4
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \n22_adj_1701_cascade_\
        );

    \I__1996\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21985\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__21985\,
            I => \N__21980\
        );

    \I__1994\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21977\
        );

    \I__1993\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21974\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__21980\,
            I => \N__21971\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21968\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__21974\,
            I => buf_adcdata_vac_7
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__21971\,
            I => buf_adcdata_vac_7
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__21968\,
            I => buf_adcdata_vac_7
        );

    \I__1987\ : InMux
    port map (
            O => \N__21961\,
            I => \N__21958\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__21958\,
            I => \N__21953\
        );

    \I__1985\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21948\
        );

    \I__1984\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21948\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__21953\,
            I => buf_adcdata_iac_4
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__21948\,
            I => buf_adcdata_iac_4
        );

    \I__1981\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21938\
        );

    \I__1980\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21935\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__21941\,
            I => \N__21932\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21929\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21926\
        );

    \I__1976\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21923\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__21929\,
            I => read_buf_14
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__21926\,
            I => read_buf_14
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__21923\,
            I => read_buf_14
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__21916\,
            I => \N__21911\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__21915\,
            I => \N__21908\
        );

    \I__1970\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21905\
        );

    \I__1969\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21902\
        );

    \I__1968\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21899\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21896\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__21902\,
            I => \N__21893\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__21899\,
            I => read_buf_3
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__21896\,
            I => read_buf_3
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__21893\,
            I => read_buf_3
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__21886\,
            I => \N__21881\
        );

    \I__1961\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21878\
        );

    \I__1960\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21873\
        );

    \I__1959\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21873\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__21878\,
            I => read_buf_13
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__21873\,
            I => read_buf_13
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__21868\,
            I => \n19_adj_1690_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21862\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__21862\,
            I => \N__21858\
        );

    \I__1953\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21854\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__21858\,
            I => \N__21851\
        );

    \I__1951\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21848\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__21854\,
            I => buf_adcdata_vac_6
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__21851\,
            I => buf_adcdata_vac_6
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__21848\,
            I => buf_adcdata_vac_6
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__21841\,
            I => \n19_adj_1693_cascade_\
        );

    \I__1946\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21833\
        );

    \I__1945\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21828\
        );

    \I__1944\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21828\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__21833\,
            I => read_buf_10
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__21828\,
            I => read_buf_10
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__21823\,
            I => \N__21819\
        );

    \I__1940\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21815\
        );

    \I__1939\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21810\
        );

    \I__1938\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21810\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21807\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__21810\,
            I => bit_cnt_2
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__21807\,
            I => bit_cnt_2
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__1933\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21793\
        );

    \I__1932\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21786\
        );

    \I__1931\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21786\
        );

    \I__1930\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21786\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21783\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__21786\,
            I => bit_cnt_1
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__21783\,
            I => bit_cnt_1
        );

    \I__1926\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21769\
        );

    \I__1925\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21769\
        );

    \I__1924\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21764\
        );

    \I__1923\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21758\
        );

    \I__1922\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21758\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21755\
        );

    \I__1920\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21751\
        );

    \I__1919\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21748\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21744\
        );

    \I__1917\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21741\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21736\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__21755\,
            I => \N__21736\
        );

    \I__1914\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21733\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__21751\,
            I => \N__21728\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__21748\,
            I => \N__21728\
        );

    \I__1911\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21725\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__21744\,
            I => dds_state_0_adj_1510
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__21741\,
            I => dds_state_0_adj_1510
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__21736\,
            I => dds_state_0_adj_1510
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__21733\,
            I => dds_state_0_adj_1510
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__21728\,
            I => dds_state_0_adj_1510
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__21725\,
            I => dds_state_0_adj_1510
        );

    \I__1904\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__21709\,
            I => n8_adj_1686
        );

    \I__1902\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21701\
        );

    \I__1901\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21698\
        );

    \I__1900\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21695\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21692\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21687\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__21695\,
            I => \N__21687\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__21692\,
            I => read_buf_11
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__21687\,
            I => read_buf_11
        );

    \I__1894\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21678\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__21681\,
            I => \N__21674\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__21678\,
            I => \N__21671\
        );

    \I__1891\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21666\
        );

    \I__1890\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21666\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__21671\,
            I => read_buf_12
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__21666\,
            I => read_buf_12
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__21661\,
            I => \RTD.n22632_cascade_\
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__21658\,
            I => \N__21655\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__1884\ : Span12Mux_s0_v
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__21649\,
            I => \DDS_CS1\
        );

    \I__1882\ : CEMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__21637\,
            I => \CLK_DDS.n9_adj_1489\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__21634\,
            I => \N__21630\
        );

    \I__1877\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21625\
        );

    \I__1876\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21625\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__21625\,
            I => read_buf_15
        );

    \I__1874\ : InMux
    port map (
            O => \N__21622\,
            I => \ADC_VAC.n20685\
        );

    \I__1873\ : InMux
    port map (
            O => \N__21619\,
            I => \ADC_VAC.n20686\
        );

    \I__1872\ : InMux
    port map (
            O => \N__21616\,
            I => \ADC_VAC.n20687\
        );

    \I__1871\ : InMux
    port map (
            O => \N__21613\,
            I => \ADC_VAC.n20688\
        );

    \I__1870\ : InMux
    port map (
            O => \N__21610\,
            I => \ADC_VAC.n20689\
        );

    \I__1869\ : CEMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__21604\,
            I => \ADC_VAC.n13784\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__21601\,
            I => \ADC_VAC.n13784_cascade_\
        );

    \I__1866\ : SRMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__21589\,
            I => \ADC_VAC.n15660\
        );

    \I__1862\ : CEMux
    port map (
            O => \N__21586\,
            I => \N__21582\
        );

    \I__1861\ : CEMux
    port map (
            O => \N__21585\,
            I => \N__21579\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__21582\,
            I => \N__21576\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__21579\,
            I => \N__21573\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__21576\,
            I => \N__21570\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__21573\,
            I => \N__21567\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__21570\,
            I => \CLK_DDS.n9\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__21567\,
            I => \CLK_DDS.n9\
        );

    \I__1854\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21559\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__21559\,
            I => \N__21556\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__21556\,
            I => \N__21551\
        );

    \I__1851\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21546\
        );

    \I__1850\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21546\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__21551\,
            I => buf_adcdata_vac_4
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__21546\,
            I => buf_adcdata_vac_4
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__1846\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21534\
        );

    \I__1845\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21531\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__21534\,
            I => cmd_rdadctmp_1_adj_1547
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__21531\,
            I => cmd_rdadctmp_1_adj_1547
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21523\
        );

    \I__1841\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__21520\,
            I => \N__21516\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__21519\,
            I => \N__21513\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__21516\,
            I => \N__21509\
        );

    \I__1837\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21504\
        );

    \I__1836\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21504\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__21509\,
            I => cmd_rdadctmp_14_adj_1534
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__21504\,
            I => cmd_rdadctmp_14_adj_1534
        );

    \I__1833\ : InMux
    port map (
            O => \N__21499\,
            I => \bfn_2_14_0_\
        );

    \I__1832\ : InMux
    port map (
            O => \N__21496\,
            I => \ADC_VAC.n20683\
        );

    \I__1831\ : InMux
    port map (
            O => \N__21493\,
            I => \ADC_VAC.n20684\
        );

    \I__1830\ : CEMux
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__21487\,
            I => \RTD.n12262\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__21484\,
            I => \N__21481\
        );

    \I__1827\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21478\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__21472\,
            I => \N__21469\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__21469\,
            I => \N__21466\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__21466\,
            I => \N__21463\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__21463\,
            I => \RTD_SDO\
        );

    \I__1820\ : SRMux
    port map (
            O => \N__21460\,
            I => \N__21457\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__21457\,
            I => \CLK_DDS.n18366\
        );

    \I__1818\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21447\
        );

    \I__1817\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21440\
        );

    \I__1816\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21440\
        );

    \I__1815\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21440\
        );

    \I__1814\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21437\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__21447\,
            I => bit_cnt_0_adj_1512
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__21440\,
            I => bit_cnt_0_adj_1512
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__21437\,
            I => bit_cnt_0_adj_1512
        );

    \I__1810\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21426\
        );

    \I__1809\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21423\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__21426\,
            I => bit_cnt_3
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__21423\,
            I => bit_cnt_3
        );

    \I__1806\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21415\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__21415\,
            I => n22326
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__1803\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21406\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21403\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__1800\ : Span4Mux_h
    port map (
            O => \N__21400\,
            I => \N__21397\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__21397\,
            I => \VAC_MISO\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__1797\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21385\
        );

    \I__1796\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21385\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__21385\,
            I => cmd_rdadctmp_0_adj_1548
        );

    \I__1794\ : IoInMux
    port map (
            O => \N__21382\,
            I => \N__21379\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21375\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__21378\,
            I => \N__21372\
        );

    \I__1791\ : Span12Mux_s4_h
    port map (
            O => \N__21375\,
            I => \N__21369\
        );

    \I__1790\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21366\
        );

    \I__1789\ : Odrv12
    port map (
            O => \N__21369\,
            I => \VAC_SCLK\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__21366\,
            I => \VAC_SCLK\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__21361\,
            I => \n14_cascade_\
        );

    \I__1786\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21355\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__21355\,
            I => n21889
        );

    \I__1784\ : IoInMux
    port map (
            O => \N__21352\,
            I => \N__21349\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__21349\,
            I => \N__21345\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__21348\,
            I => \N__21342\
        );

    \I__1781\ : Span12Mux_s4_h
    port map (
            O => \N__21345\,
            I => \N__21339\
        );

    \I__1780\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21336\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__21339\,
            I => \VAC_CS\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__21336\,
            I => \VAC_CS\
        );

    \I__1777\ : IoInMux
    port map (
            O => \N__21331\,
            I => \N__21328\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21325\
        );

    \I__1775\ : Span4Mux_s3_v
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__21322\,
            I => \N__21318\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__21318\,
            I => \N__21312\
        );

    \I__1771\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__21312\,
            I => \DDS_SCK1\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__21309\,
            I => \DDS_SCK1\
        );

    \I__1768\ : IoInMux
    port map (
            O => \N__21304\,
            I => \N__21301\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__1766\ : Span4Mux_s2_h
    port map (
            O => \N__21298\,
            I => \N__21295\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__21295\,
            I => \N__21292\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__21292\,
            I => \RTD_SCLK\
        );

    \I__1763\ : CEMux
    port map (
            O => \N__21289\,
            I => \N__21286\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__21286\,
            I => \N__21283\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__21283\,
            I => \RTD.n8\
        );

    \I__1760\ : IoInMux
    port map (
            O => \N__21280\,
            I => \N__21277\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__21277\,
            I => \N__21274\
        );

    \I__1758\ : IoSpan4Mux
    port map (
            O => \N__21274\,
            I => \N__21271\
        );

    \I__1757\ : IoSpan4Mux
    port map (
            O => \N__21271\,
            I => \N__21268\
        );

    \I__1756\ : Span4Mux_s3_h
    port map (
            O => \N__21268\,
            I => \N__21265\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__21265\,
            I => \RTD_SDI\
        );

    \I__1754\ : SRMux
    port map (
            O => \N__21262\,
            I => \N__21259\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__21259\,
            I => \RTD.n21253\
        );

    \I__1752\ : IoInMux
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__1750\ : IoSpan4Mux
    port map (
            O => \N__21250\,
            I => \N__21247\
        );

    \I__1749\ : IoSpan4Mux
    port map (
            O => \N__21247\,
            I => \N__21244\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__21244\,
            I => \ICE_SYSCLK\
        );

    \I__1747\ : IoInMux
    port map (
            O => \N__21241\,
            I => \N__21238\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__21238\,
            I => \N__21235\
        );

    \I__1745\ : IoSpan4Mux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__1744\ : Span4Mux_s3_v
    port map (
            O => \N__21232\,
            I => \N__21229\
        );

    \I__1743\ : Sp12to4
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__1742\ : Span12Mux_h
    port map (
            O => \N__21226\,
            I => \N__21223\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__21223\,
            I => \ICE_GPMO_2\
        );

    \INVADC_VDC.genclk.t0off_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i8C_net\,
            I => \N__48417\
        );

    \INVADC_VDC.genclk.t0off_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i0C_net\,
            I => \N__48416\
        );

    \INVADC_VDC.genclk.div_state_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i0C_net\,
            I => \N__48415\
        );

    \INVADC_VDC.genclk.div_state_i1C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i1C_net\,
            I => \N__48412\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__61891\
        );

    \INVdds0_mclk_297C\ : INV
    port map (
            O => \INVdds0_mclk_297C_net\,
            I => \N__48414\
        );

    \INVdds0_mclkcnt_i7_3792__i0C\ : INV
    port map (
            O => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            I => \N__48413\
        );

    \INVADC_VDC.genclk.t0on_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i8C_net\,
            I => \N__48411\
        );

    \INVADC_VDC.genclk.t0on_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i0C_net\,
            I => \N__48409\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__61973\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__61956\
        );

    \INVcomm_spi.bit_cnt_3787__i3C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_3787__i3C_net\,
            I => \N__53678\
        );

    \INVADC_VDC.genclk.t_clk_24C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t_clk_24C_net\,
            I => \N__48402\
        );

    \INVcomm_spi.MISO_48_12606_12607_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12606_12607_setC_net\,
            I => \N__61937\
        );

    \INVcomm_spi.imiso_83_12612_12613_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12612_12613_setC_net\,
            I => \N__53706\
        );

    \INVcomm_spi.MISO_48_12606_12607_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12606_12607_resetC_net\,
            I => \N__61829\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__61969\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__61951\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__61935\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__61887\
        );

    \INVeis_state_i2C\ : INV
    port map (
            O => \INVeis_state_i2C_net\,
            I => \N__61900\
        );

    \INVeis_end_302C\ : INV
    port map (
            O => \INVeis_end_302C_net\,
            I => \N__61886\
        );

    \INVcomm_spi.imiso_83_12612_12613_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12612_12613_resetC_net\,
            I => \N__53638\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__61913\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__61899\
        );

    \INVacadc_trig_303C\ : INV
    port map (
            O => \INVacadc_trig_303C_net\,
            I => \N__61947\
        );

    \INViac_raw_buf_vac_raw_buf_merged2WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            I => \N__61923\
        );

    \INViac_raw_buf_vac_raw_buf_merged7WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            I => \N__62014\
        );

    \INViac_raw_buf_vac_raw_buf_merged1WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            I => \N__61851\
        );

    \INViac_raw_buf_vac_raw_buf_merged6WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            I => \N__62011\
        );

    \INViac_raw_buf_vac_raw_buf_merged0WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            I => \N__61838\
        );

    \INViac_raw_buf_vac_raw_buf_merged5WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            I => \N__62004\
        );

    \INViac_raw_buf_vac_raw_buf_merged9WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            I => \N__61882\
        );

    \INViac_raw_buf_vac_raw_buf_merged4WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            I => \N__61989\
        );

    \INViac_raw_buf_vac_raw_buf_merged8WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            I => \N__61860\
        );

    \INViac_raw_buf_vac_raw_buf_merged10WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            I => \N__61868\
        );

    \INViac_raw_buf_vac_raw_buf_merged3WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            I => \N__61960\
        );

    \INViac_raw_buf_vac_raw_buf_merged11WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            I => \N__61893\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20773,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20781,
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20789,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20797,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20805,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n20637_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20645,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20629,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20620,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20668,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n20659,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_23_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_5_0_\
        );

    \IN_MUX_bfv_23_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n20743\,
            carryinitout => \bfn_23_6_0_\
        );

    \IN_MUX_bfv_19_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_5_0_\
        );

    \IN_MUX_bfv_19_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n20758\,
            carryinitout => \bfn_19_6_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n20732\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n20697\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n20705\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n20713\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n20721\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_16_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RTD.SCLK_51_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100000011110"
        )
    port map (
            in0 => \N__26680\,
            in1 => \N__26864\,
            in2 => \N__26521\,
            in3 => \N__26249\,
            lcout => \RTD_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35006\,
            ce => \N__21289\,
            sr => \_gnd_net_\
        );

    \RTD.i20152_4_lut_4_lut_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111011111"
        )
    port map (
            in0 => \N__26837\,
            in1 => \N__26674\,
            in2 => \N__26503\,
            in3 => \N__26223\,
            lcout => \RTD.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_4_lut_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__26866\,
            in1 => \N__26675\,
            in2 => \N__26519\,
            in3 => \N__26229\,
            lcout => \RTD.n21253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.MOSI_59_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__22657\,
            in1 => \N__26510\,
            in2 => \N__22768\,
            in3 => \N__26234\,
            lcout => \RTD_SDI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35038\,
            ce => \N__21490\,
            sr => \N__21262\
        );

    \CLK_DDS.bit_cnt_i3_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__21453\,
            in1 => \N__21798\,
            in2 => \N__21823\,
            in3 => \N__21430\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61925\,
            ce => \N__24640\,
            sr => \N__21460\
        );

    \CLK_DDS.bit_cnt_i2_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__21797\,
            in1 => \N__21452\,
            in2 => \_gnd_net_\,
            in3 => \N__21818\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61925\,
            ce => \N__24640\,
            sr => \N__21460\
        );

    \CLK_DDS.bit_cnt_i1_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21451\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21796\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61925\,
            ce => \N__24640\,
            sr => \N__21460\
        );

    \ADC_VAC.cmd_rdadctmp_i1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__21537\,
            in1 => \N__33954\,
            in2 => \N__21394\,
            in3 => \N__35925\,
            lcout => cmd_rdadctmp_1_adj_1547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__21390\,
            in1 => \N__33953\,
            in2 => \N__21412\,
            in3 => \N__35924\,
            lcout => cmd_rdadctmp_0_adj_1548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i1_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__32099\,
            in1 => \N__31992\,
            in2 => \_gnd_net_\,
            in3 => \N__35926\,
            lcout => adc_state_1_adj_1515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62009\,
            ce => \N__22267\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_303_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31970\,
            in2 => \_gnd_net_\,
            in3 => \N__32093\,
            lcout => n21889,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.SCLK_35_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011100010"
        )
    port map (
            in0 => \N__32095\,
            in1 => \N__31972\,
            in2 => \N__21378\,
            in3 => \N__35913\,
            lcout => \VAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_196_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001110"
        )
    port map (
            in0 => \N__32094\,
            in1 => \N__31971\,
            in2 => \N__21348\,
            in3 => \N__35911\,
            lcout => OPEN,
            ltout => \n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.CS_37_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__35912\,
            in1 => \N__22310\,
            in2 => \N__21361\,
            in3 => \N__21358\,
            lcout => \VAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__24704\,
            in1 => \N__21774\,
            in2 => \N__24639\,
            in3 => \N__21454\,
            lcout => bit_cnt_0_adj_1512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.SCLK_27_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011111001"
        )
    port map (
            in0 => \N__21775\,
            in1 => \N__24614\,
            in2 => \N__21321\,
            in3 => \N__24703\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i27_4_lut_4_lut_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010010100"
        )
    port map (
            in0 => \N__26862\,
            in1 => \N__26676\,
            in2 => \N__26520\,
            in3 => \N__26233\,
            lcout => \RTD.n12262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i7_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57877\,
            in1 => \N__48800\,
            in2 => \N__46654\,
            in3 => \N__35337\,
            lcout => \buf_cfgRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__22529\,
            in1 => \N__24083\,
            in2 => \N__21484\,
            in3 => \N__23976\,
            lcout => read_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i1_3_lut_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__24546\,
            in1 => \N__24691\,
            in2 => \_gnd_net_\,
            in3 => \N__21767\,
            lcout => \CLK_DDS.n18366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19900_2_lut_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21450\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21429\,
            lcout => n22326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__23975\,
            in1 => \N__22482\,
            in2 => \N__24091\,
            in3 => \N__22530\,
            lcout => read_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010100000101"
        )
    port map (
            in0 => \N__21763\,
            in1 => \N__21712\,
            in2 => \N__24609\,
            in3 => \N__21418\,
            lcout => dds_state_0_adj_1510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61926\,
            ce => \N__21585\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.i20153_4_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__24522\,
            in1 => \N__21754\,
            in2 => \N__56236\,
            in3 => \N__24706\,
            lcout => \CLK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i6_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__35946\,
            in2 => \N__21526\,
            in3 => \N__21861\,
            lcout => buf_adcdata_vac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24707\,
            in2 => \_gnd_net_\,
            in3 => \N__21768\,
            lcout => dds_state_1_adj_1509,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61961\,
            ce => \N__21586\,
            sr => \N__24635\
        );

    \ADC_VAC.ADC_DATA_i4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__21555\,
            in1 => \N__35602\,
            in2 => \N__24321\,
            in3 => \N__35923\,
            lcout => buf_adcdata_vac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61977\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_4_i19_3_lut_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24985\,
            in1 => \N__21554\,
            in2 => \_gnd_net_\,
            in3 => \N__59112\,
            lcout => n19_adj_1700,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i2_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35868\,
            in1 => \N__22698\,
            in2 => \N__21541\,
            in3 => \N__34001\,
            lcout => cmd_rdadctmp_2_adj_1546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61990\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i14_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__21512\,
            in1 => \N__33979\,
            in2 => \N__22950\,
            in3 => \N__35777\,
            lcout => cmd_rdadctmp_14_adj_1534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i15_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22205\,
            in1 => \N__33980\,
            in2 => \N__21519\,
            in3 => \N__35778\,
            lcout => cmd_rdadctmp_15_adj_1533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i13_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22943\,
            in1 => \N__33978\,
            in2 => \N__24322\,
            in3 => \N__35776\,
            lcout => cmd_rdadctmp_13_adj_1535,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.bit_cnt_i0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22375\,
            in2 => \_gnd_net_\,
            in3 => \N__21499\,
            lcout => \ADC_VAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \ADC_VAC.n20683\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i1_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22120\,
            in2 => \_gnd_net_\,
            in3 => \N__21496\,
            lcout => \ADC_VAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20683\,
            carryout => \ADC_VAC.n20684\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22132\,
            in2 => \_gnd_net_\,
            in3 => \N__21493\,
            lcout => \ADC_VAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20684\,
            carryout => \ADC_VAC.n20685\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22107\,
            in2 => \_gnd_net_\,
            in3 => \N__21622\,
            lcout => \ADC_VAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20685\,
            carryout => \ADC_VAC.n20686\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i4_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22093\,
            in2 => \_gnd_net_\,
            in3 => \N__21619\,
            lcout => \ADC_VAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20686\,
            carryout => \ADC_VAC.n20687\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i5_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22345\,
            in2 => \_gnd_net_\,
            in3 => \N__21616\,
            lcout => \ADC_VAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20687\,
            carryout => \ADC_VAC.n20688\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i6_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22387\,
            in2 => \_gnd_net_\,
            in3 => \N__21613\,
            lcout => \ADC_VAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC.n20688\,
            carryout => \ADC_VAC.n20689\,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.bit_cnt_i7_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22360\,
            in2 => \_gnd_net_\,
            in3 => \N__21610\,
            lcout => \ADC_VAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62006\,
            ce => \N__21607\,
            sr => \N__21598\
        );

    \ADC_VAC.i1_4_lut_adj_48_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010010"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__22311\,
            in2 => \N__32092\,
            in3 => \N__35715\,
            lcout => \ADC_VAC.n13784\,
            ltout => \ADC_VAC.n13784_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i12937_2_lut_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21601\,
            in3 => \N__32071\,
            lcout => \ADC_VAC.n15660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i20201_2_lut_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35716\,
            in2 => \_gnd_net_\,
            in3 => \N__22321\,
            lcout => \ADC_VAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i20130_4_lut_LC_3_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100111001100"
        )
    port map (
            in0 => \N__24610\,
            in1 => \N__24684\,
            in2 => \N__56232\,
            in3 => \N__21777\,
            lcout => \CLK_DDS.n13376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i23_4_lut_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100111"
        )
    port map (
            in0 => \N__21778\,
            in1 => \N__56228\,
            in2 => \N__24705\,
            in3 => \N__24611\,
            lcout => \CLK_DDS.n9_adj_1489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i2_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24612\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24688\,
            lcout => dds_state_2_adj_1508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i20043_3_lut_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35131\,
            in1 => \N__26654\,
            in2 => \_gnd_net_\,
            in3 => \N__32875\,
            lcout => OPEN,
            ltout => \RTD.n22632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i17362_4_lut_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__26838\,
            in2 => \N__21661\,
            in3 => \N__22429\,
            lcout => \RTD.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.CS_28_LC_3_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__24613\,
            in1 => \N__24689\,
            in2 => \_gnd_net_\,
            in3 => \N__21776\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61869\,
            ce => \N__21646\,
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i15_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21943\,
            in1 => \N__24053\,
            in2 => \N__21634\,
            in3 => \N__23979\,
            lcout => read_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i15_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__35298\,
            in1 => \N__21633\,
            in2 => \N__26518\,
            in3 => \N__23811\,
            lcout => \buf_readRTD_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i10_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21838\,
            in1 => \N__23810\,
            in2 => \N__28740\,
            in3 => \N__26486\,
            lcout => \buf_readRTD_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19153_2_lut_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26222\,
            in2 => \_gnd_net_\,
            in3 => \N__26858\,
            lcout => \RTD.n22079\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i4_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__22508\,
            in1 => \N__23980\,
            in2 => \N__21916\,
            in3 => \N__24054\,
            lcout => \RTD.read_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i10_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__21836\,
            in1 => \N__24078\,
            in2 => \N__23722\,
            in3 => \N__23982\,
            lcout => read_buf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i11_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__23981\,
            in1 => \N__21837\,
            in2 => \N__24090\,
            in3 => \N__21704\,
            lcout => read_buf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i3_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__22471\,
            in1 => \N__24079\,
            in2 => \N__21915\,
            in3 => \N__23983\,
            lcout => read_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i14_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21942\,
            in1 => \N__23816\,
            in2 => \N__23403\,
            in3 => \N__26492\,
            lcout => \buf_readRTD_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i12_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26490\,
            in1 => \N__21682\,
            in2 => \N__28851\,
            in3 => \N__23818\,
            lcout => \buf_readRTD_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i11_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21705\,
            in1 => \N__23815\,
            in2 => \N__25242\,
            in3 => \N__26491\,
            lcout => \buf_readRTD_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i3_3_lut_4_lut_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21822\,
            in1 => \N__24690\,
            in2 => \N__21802\,
            in3 => \N__21747\,
            lcout => n8_adj_1686,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i12_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21706\,
            in1 => \N__24087\,
            in2 => \N__21681\,
            in3 => \N__23985\,
            lcout => read_buf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i13_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__23984\,
            in1 => \N__21677\,
            in2 => \N__21886\,
            in3 => \N__24089\,
            lcout => read_buf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i14_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__21885\,
            in1 => \N__24088\,
            in2 => \N__21941\,
            in3 => \N__23986\,
            lcout => read_buf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i3_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26493\,
            in1 => \N__21914\,
            in2 => \N__44247\,
            in3 => \N__23817\,
            lcout => \buf_readRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i13_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21884\,
            in1 => \N__23814\,
            in2 => \N__31227\,
            in3 => \N__26494\,
            lcout => \buf_readRTD_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_7_i19_3_lut_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25027\,
            in1 => \N__21984\,
            in2 => \_gnd_net_\,
            in3 => \N__59509\,
            lcout => OPEN,
            ltout => \n19_adj_1690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_7_i22_3_lut_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22040\,
            in2 => \N__21868\,
            in3 => \N__60100\,
            lcout => n22_adj_1691,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i21_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35609\,
            in1 => \N__35865\,
            in2 => \N__23145\,
            in3 => \N__31196\,
            lcout => buf_adcdata_vac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i29_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23138\,
            in1 => \N__33902\,
            in2 => \N__23008\,
            in3 => \N__35866\,
            lcout => cmd_rdadctmp_29_adj_1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_6_i19_3_lut_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__21857\,
            in1 => \N__25183\,
            in2 => \N__59518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n19_adj_1693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_6_i22_3_lut_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22061\,
            in2 => \N__21841\,
            in3 => \N__60099\,
            lcout => n22_adj_1694,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_5_i30_3_lut_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__22081\,
            in1 => \N__22225\,
            in2 => \N__61057\,
            in3 => \_gnd_net_\,
            lcout => n30_adj_1698,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i6_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__22062\,
            in1 => \N__39406\,
            in2 => \N__22024\,
            in3 => \N__39780\,
            lcout => buf_adcdata_iac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i7_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__39775\,
            in1 => \N__22968\,
            in2 => \N__39418\,
            in3 => \N__22044\,
            lcout => buf_adcdata_iac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i14_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22019\,
            in1 => \N__39776\,
            in2 => \N__22189\,
            in3 => \N__37831\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i15_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37830\,
            in1 => \N__22020\,
            in2 => \N__39809\,
            in3 => \N__22967\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_4_i22_3_lut_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60083\,
            in1 => \N__21956\,
            in2 => \_gnd_net_\,
            in3 => \N__22009\,
            lcout => OPEN,
            ltout => \n22_adj_1701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_4_i30_3_lut_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22003\,
            in2 => \N__21991\,
            in3 => \N__61017\,
            lcout => n30_adj_1702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i7_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__35881\,
            in2 => \N__22219\,
            in3 => \N__21983\,
            lcout => buf_adcdata_vac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i4_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39386\,
            in1 => \N__39781\,
            in2 => \N__22686\,
            in3 => \N__21957\,
            lcout => buf_adcdata_iac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_5_i22_3_lut_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__22855\,
            in2 => \_gnd_net_\,
            in3 => \N__60082\,
            lcout => n22_adj_1697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i13_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22178\,
            in1 => \N__39819\,
            in2 => \N__22687\,
            in3 => \N__37832\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i16_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22808\,
            in1 => \N__35867\,
            in2 => \N__22212\,
            in3 => \N__33939\,
            lcout => cmd_rdadctmp_16_adj_1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i5_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39399\,
            in1 => \N__39818\,
            in2 => \N__22185\,
            in3 => \N__22161\,
            lcout => buf_adcdata_iac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i8_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35587\,
            in1 => \N__35775\,
            in2 => \N__22818\,
            in3 => \N__25283\,
            lcout => buf_adcdata_vac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i23_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35774\,
            in1 => \N__23040\,
            in2 => \N__24262\,
            in3 => \N__33981\,
            lcout => cmd_rdadctmp_23_adj_1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i3_3_lut_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__25876\,
            in1 => \N__32089\,
            in2 => \_gnd_net_\,
            in3 => \N__35712\,
            lcout => OPEN,
            ltout => \ADC_VAC.n13747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__31999\,
            in1 => \N__22138\,
            in2 => \N__22141\,
            in3 => \N__32090\,
            lcout => \ADC_VAC.n22030\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__22294\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35711\,
            lcout => \ADC_VAC.n13842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19182_4_lut_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22131\,
            in1 => \N__22119\,
            in2 => \N__22108\,
            in3 => \N__22092\,
            lcout => OPEN,
            ltout => \ADC_VAC.n22109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19199_4_lut_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22386\,
            in1 => \N__22374\,
            in2 => \N__22363\,
            in3 => \N__22359\,
            lcout => OPEN,
            ltout => \ADC_VAC.n22126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i20123_4_lut_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__35713\,
            in1 => \N__31991\,
            in2 => \N__22348\,
            in3 => \N__22344\,
            lcout => OPEN,
            ltout => \ADC_VAC.n22389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__32091\,
            in1 => \N__32000\,
            in2 => \N__22333\,
            in3 => \N__35714\,
            lcout => adc_state_0_adj_1516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62000\,
            ce => \N__22330\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i30_4_lut_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001101"
        )
    port map (
            in0 => \N__31998\,
            in1 => \N__22295\,
            in2 => \N__32100\,
            in3 => \N__25875\,
            lcout => \ADC_VAC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_4_lut_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000010"
        )
    port map (
            in0 => \N__31996\,
            in1 => \N__32066\,
            in2 => \N__22315\,
            in3 => \N__35709\,
            lcout => n13847,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i2_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__31997\,
            in1 => \N__32067\,
            in2 => \_gnd_net_\,
            in3 => \N__35710\,
            lcout => \DTRIG_N_1182_adj_1549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62007\,
            ce => \N__22266\,
            sr => \_gnd_net_\
        );

    \RTD.CS_52_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011111"
        )
    port map (
            in0 => \N__26672\,
            in1 => \N__22231\,
            in2 => \N__26855\,
            in3 => \N__26206\,
            lcout => \RTD_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35014\,
            ce => \N__23377\,
            sr => \_gnd_net_\
        );

    \RTD.i19756_2_lut_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23345\,
            in2 => \_gnd_net_\,
            in3 => \N__23689\,
            lcout => \RTD.n22382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_rep_43_2_lut_3_lut_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__35128\,
            in1 => \N__26646\,
            in2 => \_gnd_net_\,
            in3 => \N__32872\,
            lcout => \RTD.n23689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_21_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35129\,
            lcout => \RTD.n20051\,
            ltout => \RTD.n20051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i20050_3_lut_4_lut_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__22402\,
            in1 => \N__23202\,
            in2 => \N__22447\,
            in3 => \N__26798\,
            lcout => OPEN,
            ltout => \RTD.n22599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i3_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__22444\,
            in1 => \N__26393\,
            in2 => \N__22432\,
            in3 => \N__22428\,
            lcout => \RTD.adc_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34980\,
            ce => \N__23272\,
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i2_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__22393\,
            in1 => \N__23462\,
            in2 => \N__24940\,
            in3 => \N__26394\,
            lcout => adc_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34980\,
            ce => \N__23272\,
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_4_lut_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__32874\,
            in1 => \N__35130\,
            in2 => \N__26673\,
            in3 => \N__26799\,
            lcout => OPEN,
            ltout => \RTD.n56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100010011"
        )
    port map (
            in0 => \N__26392\,
            in1 => \N__26165\,
            in2 => \N__22414\,
            in3 => \N__22411\,
            lcout => \RTD.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34980\,
            ce => \N__23272\,
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_23_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001101"
        )
    port map (
            in0 => \N__26145\,
            in1 => \N__26785\,
            in2 => \N__26459\,
            in3 => \N__26605\,
            lcout => n13584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_26_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26604\,
            in2 => \_gnd_net_\,
            in3 => \N__26144\,
            lcout => \RTD.n71\,
            ltout => \RTD.n71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i20122_3_lut_4_lut_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__22546\,
            in1 => \N__23200\,
            in2 => \N__22396\,
            in3 => \N__26786\,
            lcout => \RTD.n22623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__26606\,
            in1 => \N__22545\,
            in2 => \N__26839\,
            in3 => \N__26146\,
            lcout => \RTD.n62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i4_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__23780\,
            in1 => \N__22515\,
            in2 => \N__30882\,
            in3 => \N__26437\,
            lcout => \buf_readRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26434\,
            in1 => \N__22537\,
            in2 => \N__25524\,
            in3 => \N__23781\,
            lcout => \buf_readRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_adj_24_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__26181\,
            in1 => \N__26433\,
            in2 => \_gnd_net_\,
            in3 => \N__26817\,
            lcout => n21989,
            ltout => \n21989_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i5_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__23939\,
            in1 => \N__22516\,
            in2 => \N__22495\,
            in3 => \N__23291\,
            lcout => read_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i2_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__24037\,
            in2 => \N__22467\,
            in3 => \N__23940\,
            lcout => read_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i1_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26435\,
            in1 => \N__22491\,
            in2 => \N__22722\,
            in3 => \N__23782\,
            lcout => \buf_readRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__23292\,
            in1 => \N__23941\,
            in2 => \N__24067\,
            in3 => \N__24107\,
            lcout => read_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26436\,
            in1 => \N__22463\,
            in2 => \N__24339\,
            in3 => \N__23783\,
            lcout => \buf_readRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__23459\,
            in1 => \N__23503\,
            in2 => \N__28965\,
            in3 => \N__22582\,
            lcout => \RTD.cfg_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i4_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__23461\,
            in2 => \N__28924\,
            in3 => \N__22591\,
            lcout => \RTD.cfg_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_20_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26185\,
            in2 => \_gnd_net_\,
            in3 => \N__26818\,
            lcout => \RTD.n68\,
            ltout => \RTD.n68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i0_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__48719\,
            in2 => \N__22594\,
            in3 => \N__22573\,
            lcout => \RTD.cfg_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_4_lut_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22590\,
            in1 => \N__22581\,
            in2 => \N__28966\,
            in3 => \N__28922\,
            lcout => \RTD.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_30_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__48720\,
            in1 => \N__22554\,
            in2 => \N__25225\,
            in3 => \N__22572\,
            lcout => OPEN,
            ltout => \RTD.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i7_4_lut_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23536\,
            in1 => \N__22564\,
            in2 => \N__22558\,
            in3 => \N__23260\,
            lcout => \RTD.adress_7_N_1009_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i3_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__23460\,
            in2 => \N__25224\,
            in3 => \N__22555\,
            lcout => \RTD.cfg_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__26670\,
            in1 => \N__26253\,
            in2 => \N__22653\,
            in3 => \N__23685\,
            lcout => \RTD.adress_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35022\,
            ce => \N__24160\,
            sr => \N__22630\
        );

    \RTD.adress_i7_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__23686\,
            in1 => \N__23598\,
            in2 => \N__26257\,
            in3 => \N__26671\,
            lcout => \RTD.adress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35022\,
            ce => \N__24160\,
            sr => \N__22630\
        );

    \RTD.i34_3_lut_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001101"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__26252\,
            in2 => \N__23363\,
            in3 => \N__23648\,
            lcout => OPEN,
            ltout => \RTD.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i35_4_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__26431\,
            in1 => \N__22624\,
            in2 => \N__22633\,
            in3 => \N__26856\,
            lcout => \RTD.n13441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19113_2_lut_3_lut_4_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__26669\,
            in1 => \N__26432\,
            in2 => \N__26248\,
            in3 => \N__26854\,
            lcout => \RTD.n15396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__26667\,
            in1 => \N__26430\,
            in2 => \_gnd_net_\,
            in3 => \N__26251\,
            lcout => \RTD.n1\,
            ltout => \RTD.n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__23649\,
            in1 => \N__23386\,
            in2 => \N__22618\,
            in3 => \N__26857\,
            lcout => \RTD.n13482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_tmp_i0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__26186\,
            in1 => \N__26499\,
            in2 => \N__48724\,
            in3 => \N__22758\,
            lcout => \RTD.cfg_tmp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__22615\,
            in1 => \N__26190\,
            in2 => \N__38245\,
            in3 => \N__26495\,
            lcout => \RTD.cfg_tmp_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i2_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__26187\,
            in1 => \N__26500\,
            in2 => \N__22609\,
            in3 => \N__28953\,
            lcout => \RTD.cfg_tmp_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__26496\,
            in1 => \N__22600\,
            in2 => \N__25217\,
            in3 => \N__26193\,
            lcout => \RTD.cfg_tmp_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i4_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__26188\,
            in1 => \N__26501\,
            in2 => \N__28923\,
            in3 => \N__22792\,
            lcout => \RTD.cfg_tmp_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__26191\,
            in2 => \N__31177\,
            in3 => \N__22786\,
            lcout => \RTD.cfg_tmp_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i6_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__26189\,
            in1 => \N__26502\,
            in2 => \N__29011\,
            in3 => \N__22780\,
            lcout => \RTD.cfg_tmp_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \RTD.cfg_tmp_i7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__26192\,
            in2 => \N__35362\,
            in3 => \N__22774\,
            lcout => \RTD.cfg_tmp_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35043\,
            ce => \N__23632\,
            sr => \N__23617\
        );

    \mux_127_Mux_6_i30_3_lut_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22747\,
            in1 => \N__22735\,
            in2 => \_gnd_net_\,
            in3 => \N__61051\,
            lcout => n30_adj_1695,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i26_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33985\,
            in1 => \N__25124\,
            in2 => \N__31551\,
            in3 => \N__35964\,
            lcout => cmd_rdadctmp_26_adj_1522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19210_3_lut_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22726\,
            in1 => \N__23842\,
            in2 => \_gnd_net_\,
            in3 => \N__60669\,
            lcout => n22137,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__33986\,
            in1 => \N__22705\,
            in2 => \N__31357\,
            in3 => \N__35965\,
            lcout => cmd_rdadctmp_3_adj_1545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i12_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__22670\,
            in2 => \N__35395\,
            in3 => \N__37801\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i19_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28805\,
            in1 => \N__33988\,
            in2 => \N__22881\,
            in3 => \N__36007\,
            lcout => cmd_rdadctmp_19_adj_1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i16_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__36003\,
            in1 => \N__35599\,
            in2 => \N__23029\,
            in3 => \N__43496\,
            lcout => buf_adcdata_vac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i10_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35598\,
            in1 => \N__36005\,
            in2 => \N__22882\,
            in3 => \N__25077\,
            lcout => buf_adcdata_vac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i9_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__36004\,
            in1 => \N__35600\,
            in2 => \N__23868\,
            in3 => \N__22896\,
            lcout => buf_adcdata_vac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_5_i19_3_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28216\,
            in1 => \N__22926\,
            in2 => \_gnd_net_\,
            in3 => \N__59111\,
            lcout => n19_adj_1696,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_7_i30_3_lut_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22846\,
            in1 => \N__22834\,
            in2 => \_gnd_net_\,
            in3 => \N__61052\,
            lcout => n30_adj_1692,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i17_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22895\,
            in1 => \N__33987\,
            in2 => \N__22822\,
            in3 => \N__36006\,
            lcout => cmd_rdadctmp_17_adj_1531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i28_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__36010\,
            in1 => \N__22994\,
            in2 => \N__27861\,
            in3 => \N__33937\,
            lcout => cmd_rdadctmp_28_adj_1520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i27_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33934\,
            in1 => \N__27854\,
            in2 => \N__25137\,
            in3 => \N__36012\,
            lcout => cmd_rdadctmp_27_adj_1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i24_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__36008\,
            in1 => \N__23021\,
            in2 => \N__23053\,
            in3 => \N__33935\,
            lcout => cmd_rdadctmp_24_adj_1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i15_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__35567\,
            in1 => \N__36011\,
            in2 => \N__24228\,
            in3 => \N__23052\,
            lcout => buf_adcdata_vac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i25_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36009\,
            in1 => \N__23022\,
            in2 => \N__31547\,
            in3 => \N__33936\,
            lcout => cmd_rdadctmp_25_adj_1523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i20_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35565\,
            in1 => \N__35922\,
            in2 => \N__23004\,
            in3 => \N__25446\,
            lcout => buf_adcdata_vac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i16_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__34589\,
            in1 => \N__39728\,
            in2 => \N__22978\,
            in3 => \N__37810\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i5_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35921\,
            in1 => \N__35566\,
            in2 => \N__22954\,
            in3 => \N__22925\,
            lcout => buf_adcdata_vac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i18_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22869\,
            in1 => \N__33950\,
            in2 => \N__22903\,
            in3 => \N__35854\,
            lcout => cmd_rdadctmp_18_adj_1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23540_bdd_4_lut_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__25411\,
            in2 => \N__32203\,
            in3 => \N__60670\,
            lcout => OPEN,
            ltout => \n23543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19349_3_lut_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23215\,
            in2 => \N__22858\,
            in3 => \N__60096\,
            lcout => n22276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i31_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23160\,
            in1 => \N__33952\,
            in2 => \N__23125\,
            in3 => \N__35917\,
            lcout => cmd_rdadctmp_31_adj_1517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i23_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__35914\,
            in1 => \N__23161\,
            in2 => \N__35571\,
            in3 => \N__23237\,
            lcout => buf_adcdata_vac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i30_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__23152\,
            in1 => \N__33951\,
            in2 => \N__23124\,
            in3 => \N__35916\,
            lcout => cmd_rdadctmp_30_adj_1518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_83_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32004\,
            in2 => \_gnd_net_\,
            in3 => \N__32072\,
            lcout => n21948,
            ltout => \n21948_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i22_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__23123\,
            in1 => \N__35915\,
            in2 => \N__23107\,
            in3 => \N__23091\,
            lcout => buf_adcdata_vac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i19_3_lut_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25162\,
            in1 => \N__23087\,
            in2 => \_gnd_net_\,
            in3 => \N__59515\,
            lcout => n19_adj_1765,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_I_0_1_lut_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39177\,
            lcout => \AC_ADC_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_4_lut_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011011000110"
        )
    port map (
            in0 => \N__26771\,
            in1 => \N__26653\,
            in2 => \N__26398\,
            in3 => \N__26174\,
            lcout => \RTD.n18274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_22_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26372\,
            in2 => \_gnd_net_\,
            in3 => \N__26117\,
            lcout => \RTD.n21988\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_2_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26608\,
            in2 => \_gnd_net_\,
            in3 => \N__23688\,
            lcout => OPEN,
            ltout => \RTD.n7_adj_1497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__23364\,
            in1 => \N__23305\,
            in2 => \N__23299\,
            in3 => \N__26791\,
            lcout => \RTD.n12274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i6_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__26375\,
            in1 => \N__43671\,
            in2 => \N__24114\,
            in3 => \N__23779\,
            lcout => \buf_readRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010000000"
        )
    port map (
            in0 => \N__26607\,
            in1 => \N__26790\,
            in2 => \N__26224\,
            in3 => \N__26373\,
            lcout => n13603,
            ltout => \n13603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i5_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__26374\,
            in1 => \N__38004\,
            in2 => \N__23296\,
            in3 => \N__23293\,
            lcout => \buf_readRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__23458\,
            in1 => \N__23515\,
            in2 => \N__26517\,
            in3 => \N__23278\,
            lcout => \RTD.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35002\,
            ce => \N__23271\,
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23526\,
            in1 => \N__23415\,
            in2 => \N__35354\,
            in3 => \N__38238\,
            lcout => \RTD.n11_adj_1500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23432_bdd_4_lut_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__23250\,
            in1 => \N__35287\,
            in2 => \N__25009\,
            in3 => \N__60649\,
            lcout => n23435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.mode_53_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__23464\,
            in1 => \N__23311\,
            in2 => \N__23201\,
            in3 => \N__23687\,
            lcout => \RTD.mode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i6_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23554\,
            in1 => \N__29009\,
            in2 => \N__23476\,
            in3 => \N__23509\,
            lcout => \RTD.cfg_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i5_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23545\,
            in1 => \N__31159\,
            in2 => \N__23474\,
            in3 => \N__23507\,
            lcout => \RTD.cfg_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_adj_29_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__23553\,
            in1 => \N__29010\,
            in2 => \N__31169\,
            in3 => \N__23544\,
            lcout => \RTD.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__23463\,
            in1 => \N__23506\,
            in2 => \N__23530\,
            in3 => \N__38237\,
            lcout => \RTD.cfg_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i17375_3_lut_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__26609\,
            in1 => \N__26863\,
            in2 => \_gnd_net_\,
            in3 => \N__26225\,
            lcout => \RTD.n20093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i7_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23416\,
            in1 => \N__23508\,
            in2 => \N__23475\,
            in3 => \N__35355\,
            lcout => \RTD.cfg_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i14786_3_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23404\,
            in1 => \N__29008\,
            in2 => \_gnd_net_\,
            in3 => \N__59246\,
            lcout => n20_adj_1766,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_28_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26473\,
            lcout => \RTD.n68_adj_1498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i20131_3_lut_3_lut_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000110100001"
        )
    port map (
            in0 => \N__26474\,
            in1 => \N__26618\,
            in2 => \N__26865\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n21954\,
            ltout => \RTD.n21954_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_4_lut_adj_31_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__23365\,
            in1 => \N__26853\,
            in2 => \N__23314\,
            in3 => \N__23650\,
            lcout => \RTD.n21955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i5_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57621\,
            in1 => \N__48810\,
            in2 => \N__45340\,
            in3 => \N__31158\,
            lcout => \buf_cfgRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_25_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26250\,
            in2 => \_gnd_net_\,
            in3 => \N__23678\,
            lcout => \RTD.n11\,
            ltout => \RTD.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i30_4_lut_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__26475\,
            in1 => \N__24946\,
            in2 => \N__23635\,
            in3 => \N__23605\,
            lcout => \RTD.n13488\,
            ltout => \RTD.n13488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12862_2_lut_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23620\,
            in3 => \N__26852\,
            lcout => \RTD.n15585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19155_2_lut_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__26848\,
            in1 => \N__26616\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n22081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i6_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__24159\,
            in1 => \N__23583\,
            in2 => \N__23599\,
            in3 => \N__24929\,
            lcout => \RTD.adress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i5_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23584\,
            in1 => \N__24924\,
            in2 => \N__23575\,
            in3 => \N__24158\,
            lcout => \RTD.adress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i4_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__24157\,
            in1 => \N__23574\,
            in2 => \N__24933\,
            in3 => \N__23563\,
            lcout => \RTD.adress_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23562\,
            in1 => \N__24923\,
            in2 => \N__24181\,
            in3 => \N__24156\,
            lcout => \RTD.adress_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__24155\,
            in1 => \N__24180\,
            in2 => \N__24133\,
            in3 => \N__24928\,
            lcout => \RTD.adress_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i9_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__23835\,
            in1 => \N__24052\,
            in2 => \N__23714\,
            in3 => \N__23974\,
            lcout => read_buf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24132\,
            in1 => \N__24922\,
            in2 => \N__24169\,
            in3 => \N__24154\,
            lcout => \RTD.adress_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i8_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__23977\,
            in1 => \N__23892\,
            in2 => \N__23836\,
            in3 => \N__24077\,
            lcout => read_buf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i7_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__24118\,
            in1 => \N__24076\,
            in2 => \N__23893\,
            in3 => \N__23978\,
            lcout => read_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i7_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__24192\,
            in1 => \N__23891\,
            in2 => \N__23812\,
            in3 => \N__26515\,
            lcout => \buf_readRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_1_i19_3_lut_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24961\,
            in1 => \N__23861\,
            in2 => \_gnd_net_\,
            in3 => \N__59466\,
            lcout => n19_adj_1752,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i8_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__26514\,
            in1 => \N__23834\,
            in2 => \N__23813\,
            in3 => \N__43305\,
            lcout => \buf_readRTD_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i9_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__38256\,
            in1 => \N__23792\,
            in2 => \N__23715\,
            in3 => \N__26516\,
            lcout => \buf_readRTD_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__35001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19222_3_lut_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__60619\,
            in1 => \N__24343\,
            in2 => \_gnd_net_\,
            in3 => \N__25051\,
            lcout => n22149,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i12_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35896\,
            in1 => \N__33669\,
            in2 => \N__34000\,
            in3 => \N__24305\,
            lcout => cmd_rdadctmp_12_adj_1536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i11_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__33668\,
            in1 => \N__33973\,
            in2 => \N__36043\,
            in3 => \N__35897\,
            lcout => cmd_rdadctmp_11_adj_1537,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i22_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24248\,
            in1 => \N__33974\,
            in2 => \N__31275\,
            in3 => \N__35898\,
            lcout => cmd_rdadctmp_22_adj_1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.MOSI_31_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24273\,
            in1 => \N__24354\,
            in2 => \_gnd_net_\,
            in3 => \N__24618\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i14_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__35909\,
            in2 => \N__24258\,
            in3 => \N__28664\,
            lcout => buf_adcdata_vac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i21_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33938\,
            in1 => \N__31268\,
            in2 => \N__28788\,
            in3 => \N__35910\,
            lcout => cmd_rdadctmp_21_adj_1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_7_i19_3_lut_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25045\,
            in1 => \N__24218\,
            in2 => \_gnd_net_\,
            in3 => \N__59475\,
            lcout => OPEN,
            ltout => \n19_adj_1714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19345_3_lut_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60665\,
            in2 => \N__24199\,
            in3 => \N__24196\,
            lcout => n22272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i10_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24619\,
            in1 => \N__24748\,
            in2 => \N__24373\,
            in3 => \N__30638\,
            lcout => \CLK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i11_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24749\,
            in1 => \N__24620\,
            in2 => \N__24415\,
            in3 => \N__29734\,
            lcout => \CLK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i12_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24621\,
            in1 => \N__24750\,
            in2 => \N__24406\,
            in3 => \N__27970\,
            lcout => \CLK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i13_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24751\,
            in1 => \N__24622\,
            in2 => \N__24397\,
            in3 => \N__55237\,
            lcout => \CLK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i14_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24623\,
            in1 => \N__24752\,
            in2 => \N__24388\,
            in3 => \N__29066\,
            lcout => \CLK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i15_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__24753\,
            in1 => \N__24624\,
            in2 => \N__25347\,
            in3 => \N__24379\,
            lcout => tmp_buf_15_adj_1511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i9_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24626\,
            in1 => \N__24755\,
            in2 => \N__24364\,
            in3 => \N__31891\,
            lcout => \CLK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i8_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24754\,
            in1 => \N__24625\,
            in2 => \N__24478\,
            in3 => \N__34150\,
            lcout => \CLK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61930\,
            ce => \N__24465\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__24628\,
            in1 => \N__24756\,
            in2 => \N__37228\,
            in3 => \N__24355\,
            lcout => \CLK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i1_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24757\,
            in1 => \N__24629\,
            in2 => \N__24817\,
            in3 => \N__42133\,
            lcout => \CLK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i2_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24630\,
            in1 => \N__24758\,
            in2 => \N__24808\,
            in3 => \N__42095\,
            lcout => \CLK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i3_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24759\,
            in1 => \N__24631\,
            in2 => \N__24799\,
            in3 => \N__36868\,
            lcout => \CLK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i4_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24632\,
            in1 => \N__24760\,
            in2 => \N__24790\,
            in3 => \N__49462\,
            lcout => \CLK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i5_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__24761\,
            in1 => \N__28722\,
            in2 => \N__24781\,
            in3 => \N__24633\,
            lcout => \CLK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i6_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__31327\,
            in1 => \N__24627\,
            in2 => \N__24772\,
            in3 => \N__24762\,
            lcout => \CLK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i7_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__24763\,
            in1 => \N__24634\,
            in2 => \N__24487\,
            in3 => \N__27908\,
            lcout => \CLK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61946\,
            ce => \N__24469\,
            sr => \_gnd_net_\
        );

    \buf_dds1_i12_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__55388\,
            in1 => \N__27968\,
            in2 => \N__44719\,
            in3 => \N__49518\,
            lcout => buf_dds1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20439_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24436\,
            in1 => \N__60098\,
            in2 => \N__24430\,
            in3 => \N__60648\,
            lcout => n23366,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i12899_2_lut_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25677\,
            in2 => \_gnd_net_\,
            in3 => \N__30425\,
            lcout => \ADC_IAC.n15622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_adj_19_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010010"
        )
    port map (
            in0 => \N__30342\,
            in1 => \N__25818\,
            in2 => \N__30432\,
            in3 => \N__39549\,
            lcout => \ADC_IAC.n13667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i2_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__39551\,
            in1 => \N__30418\,
            in2 => \_gnd_net_\,
            in3 => \N__30345\,
            lcout => \DTRIG_N_1182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61993\,
            ce => \N__25840\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i1_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__30344\,
            in1 => \_gnd_net_\,
            in2 => \N__30434\,
            in3 => \N__39552\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61993\,
            ce => \N__25840\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_61_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30410\,
            in2 => \_gnd_net_\,
            in3 => \N__30340\,
            lcout => n21892,
            ltout => \n21892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_3_lut_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25817\,
            in2 => \N__24853\,
            in3 => \N__39548\,
            lcout => n13746,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_198_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110010"
        )
    port map (
            in0 => \N__30343\,
            in1 => \N__25764\,
            in2 => \N__30433\,
            in3 => \N__39550\,
            lcout => n14_adj_1578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_74_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30411\,
            in2 => \_gnd_net_\,
            in3 => \N__30341\,
            lcout => n21951,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i0_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__39630\,
            in2 => \N__24850\,
            in3 => \N__37748\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_DDS_MCLK1_THRU_LUT4_0_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48421\,
            lcout => \GB_BUFFER_DDS_MCLK1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i8_4_lut_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__25950\,
            in1 => \N__25917\,
            in2 => \N__26884\,
            in3 => \N__26904\,
            lcout => \ADC_VDC.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i9_4_lut_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25902\,
            in1 => \N__25983\,
            in2 => \N__25969\,
            in3 => \N__25935\,
            lcout => \ADC_VDC.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12594_12595_reset_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__64557\,
            lcout => \comm_spi.n15323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53689\,
            ce => 'H',
            sr => \N__35272\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_18_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__32497\,
            in1 => \N__33582\,
            in2 => \N__33432\,
            in3 => \N__32731\,
            lcout => n13925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20024_2_lut_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33380\,
            in2 => \_gnd_net_\,
            in3 => \N__32732\,
            lcout => n22388,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.SCLK_46_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__24886\,
            in1 => \N__24864\,
            in2 => \N__24895\,
            in3 => \N__32505\,
            lcout => \VDC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i12_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__27054\,
            in1 => \N__28391\,
            in2 => \N__27502\,
            in3 => \N__32723\,
            lcout => cmd_rdadctmp_12_adj_1562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i7_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__32722\,
            in1 => \N__27129\,
            in2 => \N__28401\,
            in3 => \N__27159\,
            lcout => cmd_rdadctmp_7_adj_1567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i11_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__27053\,
            in1 => \N__27084\,
            in2 => \N__32733\,
            in3 => \N__28390\,
            lcout => cmd_rdadctmp_11_adj_1563,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i2_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28386\,
            in1 => \N__32715\,
            in2 => \N__27007\,
            in3 => \N__26970\,
            lcout => cmd_rdadctmp_2_adj_1572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i8_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__27128\,
            in1 => \N__28421\,
            in2 => \N__32734\,
            in3 => \N__28392\,
            lcout => cmd_rdadctmp_8_adj_1566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28385\,
            in1 => \N__32714\,
            in2 => \N__27006\,
            in3 => \N__27033\,
            lcout => cmd_rdadctmp_1_adj_1573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i14_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27459\,
            in1 => \N__27437\,
            in2 => \N__28394\,
            in3 => \N__32712\,
            lcout => cmd_rdadctmp_14_adj_1560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31083\,
            in1 => \N__33436\,
            in2 => \N__33627\,
            in3 => \N__27475\,
            lcout => buf_adcdata_vdc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i16_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__27359\,
            in1 => \N__27412\,
            in2 => \N__28395\,
            in3 => \N__32713\,
            lcout => cmd_rdadctmp_16_adj_1558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i21_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32710\,
            in1 => \N__28372\,
            in2 => \N__27601\,
            in3 => \N__27636\,
            lcout => cmd_rdadctmp_21_adj_1553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i10_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__27083\,
            in1 => \N__28285\,
            in2 => \N__28393\,
            in3 => \N__32711\,
            lcout => cmd_rdadctmp_10_adj_1564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i13_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32708\,
            in1 => \N__27458\,
            in2 => \N__27501\,
            in3 => \N__28370\,
            lcout => cmd_rdadctmp_13_adj_1561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i20132_4_lut_4_lut_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100001"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__33586\,
            in2 => \N__33448\,
            in3 => \N__32707\,
            lcout => n12356,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i20_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32709\,
            in1 => \N__27635\,
            in2 => \N__27262\,
            in3 => \N__28371\,
            lcout => cmd_rdadctmp_20_adj_1554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i22_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32725\,
            in1 => \N__28380\,
            in2 => \N__30795\,
            in3 => \N__27599\,
            lcout => cmd_rdadctmp_22_adj_1552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i31_3_lut_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26846\,
            in1 => \N__26650\,
            in2 => \_gnd_net_\,
            in3 => \N__26235\,
            lcout => \RTD.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26847\,
            lcout => \RTD.n79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i18_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32724\,
            in1 => \N__27294\,
            in2 => \N__27337\,
            in3 => \N__28379\,
            lcout => cmd_rdadctmp_18_adj_1556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i17_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__27332\,
            in1 => \N__27360\,
            in2 => \N__28396\,
            in3 => \N__32726\,
            lcout => cmd_rdadctmp_17_adj_1557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i19_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27293\,
            in1 => \N__27260\,
            in2 => \N__28397\,
            in3 => \N__32727\,
            lcout => cmd_rdadctmp_19_adj_1555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i12_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31074\,
            in1 => \N__33443\,
            in2 => \N__30945\,
            in3 => \N__27553\,
            lcout => buf_adcdata_vdc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i17_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33440\,
            in1 => \N__31078\,
            in2 => \N__48561\,
            in3 => \N__27718\,
            lcout => buf_adcdata_vdc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i15_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31076\,
            in1 => \N__33445\,
            in2 => \N__25044\,
            in3 => \N__27520\,
            lcout => buf_adcdata_vdc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i19_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33441\,
            in1 => \N__31079\,
            in2 => \N__27753\,
            in3 => \N__27688\,
            lcout => buf_adcdata_vdc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i7_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31077\,
            in1 => \N__33446\,
            in2 => \N__25026\,
            in3 => \N__27277\,
            lcout => buf_adcdata_vdc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i23_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33442\,
            in1 => \N__31080\,
            in2 => \N__25002\,
            in3 => \N__28474\,
            lcout => buf_adcdata_vdc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i14_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31075\,
            in1 => \N__33444\,
            in2 => \N__28692\,
            in3 => \N__27535\,
            lcout => buf_adcdata_vdc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i4_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__27379\,
            in1 => \N__31081\,
            in2 => \N__24978\,
            in3 => \N__33447\,
            lcout => buf_adcdata_vdc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i10_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33394\,
            in1 => \N__31066\,
            in2 => \N__25104\,
            in3 => \N__27577\,
            lcout => buf_adcdata_vdc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i18_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33395\,
            in1 => \N__31067\,
            in2 => \N__31512\,
            in3 => \N__27703\,
            lcout => buf_adcdata_vdc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i9_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27619\,
            in1 => \N__24957\,
            in2 => \N__31084\,
            in3 => \N__33402\,
            lcout => buf_adcdata_vdc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i8_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__27238\,
            in1 => \N__25311\,
            in2 => \N__33437\,
            in3 => \N__31072\,
            lcout => buf_adcdata_vdc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i6_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31065\,
            in1 => \N__33398\,
            in2 => \N__25179\,
            in3 => \N__27313\,
            lcout => buf_adcdata_vdc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i22_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33396\,
            in1 => \N__31068\,
            in2 => \N__25158\,
            in3 => \N__27655\,
            lcout => buf_adcdata_vdc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i20_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31064\,
            in1 => \N__33397\,
            in2 => \N__25476\,
            in3 => \N__27673\,
            lcout => buf_adcdata_vdc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i18_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35992\,
            in1 => \N__35597\,
            in2 => \N__25141\,
            in3 => \N__31484\,
            lcout => buf_adcdata_vac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i112_3_lut_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60543\,
            in1 => \N__34098\,
            in2 => \_gnd_net_\,
            in3 => \N__31405\,
            lcout => OPEN,
            ltout => \n112_adj_1786_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i127_3_lut_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61412\,
            in2 => \N__25108\,
            in3 => \N__27802\,
            lcout => \comm_buf_0_7_N_543_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i11_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35596\,
            in1 => \N__35993\,
            in2 => \N__28821\,
            in3 => \N__41208\,
            lcout => buf_adcdata_vac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_2_i19_3_lut_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__25076\,
            in2 => \_gnd_net_\,
            in3 => \N__59335\,
            lcout => n19_adj_1747,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i111_3_lut_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59336\,
            in1 => \N__25356\,
            in2 => \_gnd_net_\,
            in3 => \N__34321\,
            lcout => n111_adj_1771,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i22_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__25357\,
            in1 => \N__40526\,
            in2 => \N__57869\,
            in3 => \N__45422\,
            lcout => comm_test_buf_24_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i12_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35608\,
            in1 => \N__36013\,
            in2 => \N__28789\,
            in3 => \N__30911\,
            lcout => buf_adcdata_vac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i15_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__49561\,
            in1 => \N__25340\,
            in2 => \N__46662\,
            in3 => \N__55432\,
            lcout => buf_dds1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i112_3_lut_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34299\,
            in1 => \N__60615\,
            in2 => \_gnd_net_\,
            in3 => \N__25321\,
            lcout => n112_adj_1772,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__56850\,
            in1 => \N__48814\,
            in2 => \_gnd_net_\,
            in3 => \N__25197\,
            lcout => \buf_cfgRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i14_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__29067\,
            in1 => \N__55371\,
            in2 => \N__40570\,
            in3 => \N__49560\,
            lcout => buf_dds1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_0_i19_3_lut_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25315\,
            in1 => \N__25290\,
            in2 => \_gnd_net_\,
            in3 => \N__59467\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_6_i127_3_lut_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34300\,
            in1 => \N__25261\,
            in2 => \_gnd_net_\,
            in3 => \N__61394\,
            lcout => \comm_buf_2_7_N_575_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i20_3_lut_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25249\,
            in1 => \N__25196\,
            in2 => \_gnd_net_\,
            in3 => \N__59468\,
            lcout => n20_adj_1790,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20543_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__27736\,
            in1 => \N__60080\,
            in2 => \N__25489\,
            in3 => \N__60611\,
            lcout => OPEN,
            ltout => \n23498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23498_bdd_4_lut_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__60081\,
            in1 => \N__25423\,
            in2 => \N__25480\,
            in3 => \N__25417\,
            lcout => n23501,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i19_3_lut_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59490\,
            in1 => \N__25477\,
            in2 => \_gnd_net_\,
            in3 => \N__25445\,
            lcout => n19_adj_1780,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i16_3_lut_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59488\,
            in1 => \N__29733\,
            in2 => \_gnd_net_\,
            in3 => \N__32903\,
            lcout => n16_adj_1787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i17_3_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27993\,
            in1 => \N__29799\,
            in2 => \_gnd_net_\,
            in3 => \N__59489\,
            lcout => n17_adj_1788,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__59491\,
            in1 => \N__31602\,
            in2 => \N__25392\,
            in3 => \N__60610\,
            lcout => n23540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i10_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__49567\,
            in1 => \N__30639\,
            in2 => \N__40947\,
            in3 => \N__55369\,
            lcout => buf_dds1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i23_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39351\,
            in1 => \N__39651\,
            in2 => \N__25372\,
            in3 => \N__25388\,
            lcout => buf_adcdata_iac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i7_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__55368\,
            in1 => \N__27909\,
            in2 => \N__55849\,
            in3 => \N__49569\,
            lcout => buf_dds1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i31_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__31797\,
            in1 => \N__39652\,
            in2 => \N__25371\,
            in3 => \N__37772\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20377_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25543\,
            in1 => \N__60076\,
            in2 => \N__25534\,
            in3 => \N__60609\,
            lcout => n23300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i2_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__49568\,
            in1 => \N__42096\,
            in2 => \N__52935\,
            in3 => \N__55370\,
            lcout => buf_dds1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19116_4_lut_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__45809\,
            in1 => \N__34700\,
            in2 => \N__34798\,
            in3 => \N__39170\,
            lcout => OPEN,
            ltout => \n22041_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_303_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__34701\,
            in1 => \N__45810\,
            in2 => \N__25507\,
            in3 => \N__25867\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_303C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.bit_cnt_i0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25585\,
            in2 => \_gnd_net_\,
            in3 => \N__25504\,
            lcout => \ADC_IAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \ADC_IAC.n20676\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25623\,
            in2 => \_gnd_net_\,
            in3 => \N__25501\,
            lcout => \ADC_IAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20676\,
            carryout => \ADC_IAC.n20677\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25609\,
            in2 => \_gnd_net_\,
            in3 => \N__25498\,
            lcout => \ADC_IAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20677\,
            carryout => \ADC_IAC.n20678\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25636\,
            in2 => \_gnd_net_\,
            in3 => \N__25495\,
            lcout => \ADC_IAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20678\,
            carryout => \ADC_IAC.n20679\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i4_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25648\,
            in2 => \_gnd_net_\,
            in3 => \N__25492\,
            lcout => \ADC_IAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20679\,
            carryout => \ADC_IAC.n20680\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25558\,
            in2 => \_gnd_net_\,
            in3 => \N__25696\,
            lcout => \ADC_IAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20680\,
            carryout => \ADC_IAC.n20681\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i6_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25597\,
            in2 => \_gnd_net_\,
            in3 => \N__25693\,
            lcout => \ADC_IAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_IAC.n20681\,
            carryout => \ADC_IAC.n20682\,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.bit_cnt_i7_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25570\,
            in2 => \_gnd_net_\,
            in3 => \N__25690\,
            lcout => \ADC_IAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61965\,
            ce => \N__25687\,
            sr => \N__25666\
        );

    \ADC_IAC.i1_2_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25654\,
            lcout => \ADC_IAC.n22032\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__39553\,
            in2 => \N__25819\,
            in3 => \N__25868\,
            lcout => \ADC_IAC.n22031\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19186_4_lut_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25647\,
            in1 => \N__25635\,
            in2 => \N__25624\,
            in3 => \N__25608\,
            lcout => OPEN,
            ltout => \ADC_IAC.n22113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19201_4_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25596\,
            in1 => \N__25584\,
            in2 => \N__25573\,
            in3 => \N__25569\,
            lcout => OPEN,
            ltout => \ADC_IAC.n22128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19757_4_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__39555\,
            in1 => \N__25557\,
            in2 => \N__25546\,
            in3 => \N__30367\,
            lcout => OPEN,
            ltout => \ADC_IAC.n22384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i0_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__30424\,
            in1 => \N__30366\,
            in2 => \N__25888\,
            in3 => \N__39556\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61980\,
            ce => \N__25885\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.i30_4_lut_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110000001"
        )
    port map (
            in0 => \N__25869\,
            in1 => \N__30423\,
            in2 => \N__30372\,
            in3 => \N__25816\,
            lcout => OPEN,
            ltout => \ADC_IAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i20195_2_lut_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25843\,
            in3 => \N__39554\,
            lcout => \ADC_IAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.CS_37_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__25831\,
            in1 => \N__25825\,
            in2 => \N__39715\,
            in3 => \N__25812\,
            lcout => \IAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i2_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25752\,
            in1 => \N__39622\,
            in2 => \N__25708\,
            in3 => \N__37746\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37743\,
            in1 => \N__25743\,
            in2 => \N__39713\,
            in3 => \N__25753\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__25744\,
            in1 => \N__39623\,
            in2 => \N__25735\,
            in3 => \N__37747\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37744\,
            in1 => \N__30480\,
            in2 => \N__39714\,
            in3 => \N__25734\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i1_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25704\,
            in1 => \N__39621\,
            in2 => \N__25723\,
            in3 => \N__37745\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \EIS_SYNCCLK_I_0_1_lut_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \IAC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.avg_cnt_i0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28045\,
            in2 => \_gnd_net_\,
            in3 => \N__25987\,
            lcout => \ADC_VDC.avg_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \ADC_VDC.n20725\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25984\,
            in2 => \_gnd_net_\,
            in3 => \N__25972\,
            lcout => \ADC_VDC.avg_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20725\,
            carryout => \ADC_VDC.n20726\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i2_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25968\,
            in2 => \_gnd_net_\,
            in3 => \N__25954\,
            lcout => \ADC_VDC.avg_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20726\,
            carryout => \ADC_VDC.n20727\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i3_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25951\,
            in2 => \_gnd_net_\,
            in3 => \N__25939\,
            lcout => \ADC_VDC.avg_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20727\,
            carryout => \ADC_VDC.n20728\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i4_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25936\,
            in2 => \_gnd_net_\,
            in3 => \N__25924\,
            lcout => \ADC_VDC.avg_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20728\,
            carryout => \ADC_VDC.n20729\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i5_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28033\,
            in2 => \_gnd_net_\,
            in3 => \N__25921\,
            lcout => \ADC_VDC.avg_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20729\,
            carryout => \ADC_VDC.n20730\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i6_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25918\,
            in2 => \_gnd_net_\,
            in3 => \N__25906\,
            lcout => \ADC_VDC.avg_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20730\,
            carryout => \ADC_VDC.n20731\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i7_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25903\,
            in2 => \_gnd_net_\,
            in3 => \N__25891\,
            lcout => \ADC_VDC.avg_cnt_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20731\,
            carryout => \ADC_VDC.n20732\,
            clk => \N__42747\,
            ce => \N__28637\,
            sr => \N__28563\
        );

    \ADC_VDC.avg_cnt_i8_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28017\,
            in2 => \_gnd_net_\,
            in3 => \N__26908\,
            lcout => \ADC_VDC.avg_cnt_8\,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \ADC_VDC.n20733\,
            clk => \N__42737\,
            ce => \N__28636\,
            sr => \N__28562\
        );

    \ADC_VDC.avg_cnt_i9_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26905\,
            in2 => \_gnd_net_\,
            in3 => \N__26893\,
            lcout => \ADC_VDC.avg_cnt_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20733\,
            carryout => \ADC_VDC.n20734\,
            clk => \N__42737\,
            ce => \N__28636\,
            sr => \N__28562\
        );

    \ADC_VDC.avg_cnt_i10_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28180\,
            in2 => \_gnd_net_\,
            in3 => \N__26890\,
            lcout => \ADC_VDC.avg_cnt_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20734\,
            carryout => \ADC_VDC.n20735\,
            clk => \N__42737\,
            ce => \N__28636\,
            sr => \N__28562\
        );

    \ADC_VDC.avg_cnt_i11_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26880\,
            in2 => \_gnd_net_\,
            in3 => \N__26887\,
            lcout => \ADC_VDC.avg_cnt_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42737\,
            ce => \N__28636\,
            sr => \N__28562\
        );

    \ADC_VDC.i1_4_lut_4_lut_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110010"
        )
    port map (
            in0 => \N__32607\,
            in1 => \N__28123\,
            in2 => \N__33381\,
            in3 => \N__30673\,
            lcout => \ADC_VDC.n13865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_27_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000110"
        )
    port map (
            in0 => \N__26822\,
            in1 => \N__26652\,
            in2 => \N__26472\,
            in3 => \N__26213\,
            lcout => \RTD.n18275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19145_2_lut_3_lut_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32828\,
            in1 => \N__32486\,
            in2 => \_gnd_net_\,
            in3 => \N__33516\,
            lcout => \ADC_VDC.n22071\,
            ltout => \ADC_VDC.n22071_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i34_3_lut_4_lut_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__32606\,
            in1 => \N__33552\,
            in2 => \N__26041\,
            in3 => \N__32829\,
            lcout => \ADC_VDC.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i4_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32619\,
            in1 => \N__27218\,
            in2 => \N__26941\,
            in3 => \N__28344\,
            lcout => cmd_rdadctmp_4_adj_1570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__27219\,
            in1 => \N__27188\,
            in2 => \N__28381\,
            in3 => \N__32622\,
            lcout => cmd_rdadctmp_5_adj_1569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__27439\,
            in2 => \N__27410\,
            in3 => \N__28342\,
            lcout => cmd_rdadctmp_15_adj_1559,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__32620\,
            in1 => \N__28338\,
            in2 => \N__27193\,
            in3 => \N__27158\,
            lcout => cmd_rdadctmp_6_adj_1568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__28337\,
            in1 => \N__27032\,
            in2 => \N__32800\,
            in3 => \N__32621\,
            lcout => cmd_rdadctmp_0_adj_1574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i3_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__32618\,
            in1 => \N__26969\,
            in2 => \N__26940\,
            in3 => \N__28343\,
            lcout => cmd_rdadctmp_3_adj_1571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27013\,
            in2 => \N__27034\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.cmd_rdadcbuf_0\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \ADC_VDC.n20690\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26983\,
            in2 => \N__27005\,
            in3 => \N__26977\,
            lcout => \ADC_VDC.cmd_rdadcbuf_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20690\,
            carryout => \ADC_VDC.n20691\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26950\,
            in2 => \N__26974\,
            in3 => \N__26944\,
            lcout => \ADC_VDC.cmd_rdadcbuf_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20691\,
            carryout => \ADC_VDC.n20692\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26917\,
            in2 => \N__26939\,
            in3 => \N__26911\,
            lcout => \ADC_VDC.cmd_rdadcbuf_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20692\,
            carryout => \ADC_VDC.n20693\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27202\,
            in2 => \N__27220\,
            in3 => \N__27196\,
            lcout => \ADC_VDC.cmd_rdadcbuf_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20693\,
            carryout => \ADC_VDC.n20694\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27172\,
            in2 => \N__27192\,
            in3 => \N__27163\,
            lcout => \ADC_VDC.cmd_rdadcbuf_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20694\,
            carryout => \ADC_VDC.n20695\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27139\,
            in2 => \N__27160\,
            in3 => \N__27133\,
            lcout => \ADC_VDC.cmd_rdadcbuf_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20695\,
            carryout => \ADC_VDC.n20696\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27112\,
            in2 => \N__27130\,
            in3 => \N__27106\,
            lcout => \ADC_VDC.cmd_rdadcbuf_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20696\,
            carryout => \ADC_VDC.n20697\,
            clk => \N__42738\,
            ce => \N__28626\,
            sr => \N__28557\
        );

    \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27103\,
            in2 => \N__28425\,
            in3 => \N__27097\,
            lcout => \ADC_VDC.cmd_rdadcbuf_8\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \ADC_VDC.n20698\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27094\,
            in2 => \N__28281\,
            in3 => \N__27088\,
            lcout => \ADC_VDC.cmd_rdadcbuf_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20698\,
            carryout => \ADC_VDC.n20699\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27064\,
            in2 => \N__27085\,
            in3 => \N__27058\,
            lcout => \ADC_VDC.cmd_rdadcbuf_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20699\,
            carryout => \ADC_VDC.n20700\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30957\,
            in2 => \N__27055\,
            in3 => \N__27037\,
            lcout => cmd_rdadcbuf_11,
            ltout => OPEN,
            carryin => \ADC_VDC.n20700\,
            carryout => \ADC_VDC.n20701\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27474\,
            in2 => \N__27500\,
            in3 => \N__27463\,
            lcout => cmd_rdadcbuf_12,
            ltout => OPEN,
            carryin => \ADC_VDC.n20701\,
            carryout => \ADC_VDC.n20702\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28242\,
            in2 => \N__27460\,
            in3 => \N__27442\,
            lcout => cmd_rdadcbuf_13,
            ltout => OPEN,
            carryin => \ADC_VDC.n20702\,
            carryout => \ADC_VDC.n20703\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28437\,
            in2 => \N__27438\,
            in3 => \N__27415\,
            lcout => cmd_rdadcbuf_14,
            ltout => OPEN,
            carryin => \ADC_VDC.n20703\,
            carryout => \ADC_VDC.n20704\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27375\,
            in2 => \N__27411\,
            in3 => \N__27364\,
            lcout => cmd_rdadcbuf_15,
            ltout => OPEN,
            carryin => \ADC_VDC.n20704\,
            carryout => \ADC_VDC.n20705\,
            clk => \N__42718\,
            ce => \N__28625\,
            sr => \N__28553\
        );

    \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28227\,
            in2 => \N__27361\,
            in3 => \N__27340\,
            lcout => cmd_rdadcbuf_16,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \ADC_VDC.n20706\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27309\,
            in2 => \N__27336\,
            in3 => \N__27298\,
            lcout => cmd_rdadcbuf_17,
            ltout => OPEN,
            carryin => \ADC_VDC.n20706\,
            carryout => \ADC_VDC.n20707\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27276\,
            in2 => \N__27295\,
            in3 => \N__27265\,
            lcout => cmd_rdadcbuf_18,
            ltout => OPEN,
            carryin => \ADC_VDC.n20707\,
            carryout => \ADC_VDC.n20708\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27234\,
            in2 => \N__27261\,
            in3 => \N__27223\,
            lcout => cmd_rdadcbuf_19,
            ltout => OPEN,
            carryin => \ADC_VDC.n20708\,
            carryout => \ADC_VDC.n20709\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27615\,
            in2 => \N__27637\,
            in3 => \N__27604\,
            lcout => cmd_rdadcbuf_20,
            ltout => OPEN,
            carryin => \ADC_VDC.n20709\,
            carryout => \ADC_VDC.n20710\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27576\,
            in2 => \N__27600\,
            in3 => \N__27559\,
            lcout => cmd_rdadcbuf_21,
            ltout => OPEN,
            carryin => \ADC_VDC.n20710\,
            carryout => \ADC_VDC.n20711\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28254\,
            in2 => \N__30794\,
            in3 => \N__27556\,
            lcout => cmd_rdadcbuf_22,
            ltout => OPEN,
            carryin => \ADC_VDC.n20711\,
            carryout => \ADC_VDC.n20712\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27552\,
            in2 => \N__30760\,
            in3 => \N__27541\,
            lcout => cmd_rdadcbuf_23,
            ltout => OPEN,
            carryin => \ADC_VDC.n20712\,
            carryout => \ADC_VDC.n20713\,
            clk => \N__42740\,
            ce => \N__28638\,
            sr => \N__28549\
        );

    \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31095\,
            in2 => \_gnd_net_\,
            in3 => \N__27538\,
            lcout => cmd_rdadcbuf_24,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \ADC_VDC.n20714\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27534\,
            in2 => \_gnd_net_\,
            in3 => \N__27523\,
            lcout => cmd_rdadcbuf_25,
            ltout => OPEN,
            carryin => \ADC_VDC.n20714\,
            carryout => \ADC_VDC.n20715\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27519\,
            in2 => \_gnd_net_\,
            in3 => \N__27508\,
            lcout => cmd_rdadcbuf_26,
            ltout => OPEN,
            carryin => \ADC_VDC.n20715\,
            carryout => \ADC_VDC.n20716\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28191\,
            in2 => \_gnd_net_\,
            in3 => \N__27505\,
            lcout => cmd_rdadcbuf_27,
            ltout => OPEN,
            carryin => \ADC_VDC.n20716\,
            carryout => \ADC_VDC.n20717\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27717\,
            in2 => \_gnd_net_\,
            in3 => \N__27706\,
            lcout => cmd_rdadcbuf_28,
            ltout => OPEN,
            carryin => \ADC_VDC.n20717\,
            carryout => \ADC_VDC.n20718\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__27691\,
            lcout => cmd_rdadcbuf_29,
            ltout => OPEN,
            carryin => \ADC_VDC.n20718\,
            carryout => \ADC_VDC.n20719\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27687\,
            in2 => \_gnd_net_\,
            in3 => \N__27676\,
            lcout => cmd_rdadcbuf_30,
            ltout => OPEN,
            carryin => \ADC_VDC.n20719\,
            carryout => \ADC_VDC.n20720\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27672\,
            in2 => \_gnd_net_\,
            in3 => \N__27661\,
            lcout => cmd_rdadcbuf_31,
            ltout => OPEN,
            carryin => \ADC_VDC.n20720\,
            carryout => \ADC_VDC.n20721\,
            clk => \N__42720\,
            ce => \N__28621\,
            sr => \N__28561\
        );

    \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31125\,
            in2 => \_gnd_net_\,
            in3 => \N__27658\,
            lcout => cmd_rdadcbuf_32,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \ADC_VDC.n20722\,
            clk => \N__42758\,
            ce => \N__28642\,
            sr => \N__28564\
        );

    \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27654\,
            in2 => \_gnd_net_\,
            in3 => \N__27643\,
            lcout => cmd_rdadcbuf_33,
            ltout => OPEN,
            carryin => \ADC_VDC.n20722\,
            carryout => \ADC_VDC.n20723\,
            clk => \N__42758\,
            ce => \N__28642\,
            sr => \N__28564\
        );

    \ADC_VDC.add_23_36_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28466\,
            in2 => \_gnd_net_\,
            in3 => \N__27640\,
            lcout => \ADC_VDC.cmd_rdadcbuf_35_N_1344_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12640_12641_reset_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36615\,
            in1 => \N__36591\,
            in2 => \_gnd_net_\,
            in3 => \N__36564\,
            lcout => \comm_spi.n15369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53665\,
            ce => 'H',
            sr => \N__34114\
        );

    \comm_cmd_1__bdd_4_lut_20533_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__60642\,
            in1 => \N__49705\,
            in2 => \N__60091\,
            in3 => \N__53026\,
            lcout => OPEN,
            ltout => \n23474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23474_bdd_4_lut_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__39835\,
            in1 => \N__27763\,
            in2 => \N__27808\,
            in3 => \N__60052\,
            lcout => OPEN,
            ltout => \n23477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1662065_i1_3_lut_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27724\,
            in2 => \N__27805\,
            in3 => \N__61053\,
            lcout => n30_adj_1784,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1662668_i1_3_lut_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__61054\,
            in1 => \N__29032\,
            in2 => \_gnd_net_\,
            in3 => \N__28756\,
            lcout => OPEN,
            ltout => \n30_adj_1768_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i127_3_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__61390\,
            in1 => \N__27796\,
            in2 => \N__27787\,
            in3 => \_gnd_net_\,
            lcout => \comm_buf_0_7_N_543_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20483_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__27784\,
            in1 => \N__60048\,
            in2 => \N__28834\,
            in3 => \N__60641\,
            lcout => n23426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_4_i127_3_lut_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__34102\,
            in1 => \N__27778\,
            in2 => \N__61413\,
            in3 => \_gnd_net_\,
            lcout => \comm_buf_2_7_N_575_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20034_2_lut_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59350\,
            in2 => \_gnd_net_\,
            in3 => \N__38698\,
            lcout => n22358,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i19_3_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27824\,
            in1 => \N__27757\,
            in2 => \_gnd_net_\,
            in3 => \N__59483\,
            lcout => n19_adj_1789,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23426_bdd_4_lut_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__27730\,
            in1 => \N__36814\,
            in2 => \N__27946\,
            in3 => \N__60094\,
            lcout => n23429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_337_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__59484\,
            in1 => \N__52927\,
            in2 => \N__40978\,
            in3 => \N__37403\,
            lcout => n11983,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i9_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__31877\,
            in1 => \N__55431\,
            in2 => \N__44646\,
            in3 => \N__49562\,
            lcout => buf_dds1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i11_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32904\,
            in1 => \N__56854\,
            in2 => \_gnd_net_\,
            in3 => \N__50753\,
            lcout => buf_dds0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i27_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30287\,
            in1 => \N__39754\,
            in2 => \N__27934\,
            in3 => \N__37814\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i5_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__28718\,
            in1 => \N__55403\,
            in2 => \N__47113\,
            in3 => \N__63783\,
            lcout => buf_dds1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i14_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57870\,
            in1 => \N__50764\,
            in2 => \N__40564\,
            in3 => \N__32231\,
            lcout => buf_dds0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i19_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35988\,
            in1 => \N__35603\,
            in2 => \N__27868\,
            in3 => \N__27828\,
            lcout => buf_adcdata_vac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__55402\,
            in1 => \N__37220\,
            in2 => \N__49150\,
            in3 => \N__49563\,
            lcout => buf_dds1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i13_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39341\,
            in1 => \N__39753\,
            in2 => \N__28096\,
            in3 => \N__52319\,
            lcout => buf_adcdata_iac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i6_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47077\,
            in1 => \N__50763\,
            in2 => \_gnd_net_\,
            in3 => \N__31829\,
            lcout => buf_dds0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i1_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__42125\,
            in1 => \N__55423\,
            in2 => \N__52134\,
            in3 => \N__49570\,
            lcout => buf_dds1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i19_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39402\,
            in1 => \N__39745\,
            in2 => \N__30303\,
            in3 => \N__27992\,
            lcout => buf_adcdata_iac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i16_3_lut_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32283\,
            in1 => \N__27969\,
            in2 => \_gnd_net_\,
            in3 => \N__59492\,
            lcout => n16_adj_1778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i22_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39403\,
            in1 => \N__39746\,
            in2 => \N__31801\,
            in3 => \N__31676\,
            lcout => buf_adcdata_iac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i14_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39360\,
            in1 => \N__39618\,
            in2 => \N__41297\,
            in3 => \N__28075\,
            lcout => buf_adcdata_iac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i18_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39617\,
            in1 => \N__39361\,
            in2 => \N__30603\,
            in3 => \N__27927\,
            lcout => buf_adcdata_iac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i26_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27926\,
            in1 => \N__39619\,
            in2 => \N__30460\,
            in3 => \N__37815\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_7_i16_3_lut_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27913\,
            in1 => \N__32314\,
            in2 => \_gnd_net_\,
            in3 => \N__59516\,
            lcout => n16_adj_1713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.SCLK_35_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__39608\,
            in1 => \N__30436\,
            in2 => \N__27885\,
            in3 => \N__30371\,
            lcout => \IAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i23_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37790\,
            in1 => \N__28055\,
            in2 => \N__39712\,
            in3 => \N__28074\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i21_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__28088\,
            in1 => \N__39609\,
            in2 => \N__37258\,
            in3 => \N__37791\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i22_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37789\,
            in1 => \N__28073\,
            in2 => \N__39711\,
            in3 => \N__28089\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i24_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30506\,
            in1 => \N__39610\,
            in2 => \N__28060\,
            in3 => \N__37792\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i15_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39334\,
            in1 => \N__39620\,
            in2 => \N__46910\,
            in3 => \N__28059\,
            lcout => buf_adcdata_iac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i18_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29750\,
            in1 => \N__39632\,
            in2 => \N__39216\,
            in3 => \N__37823\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i25_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37821\,
            in1 => \N__30452\,
            in2 => \N__30511\,
            in3 => \N__39636\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i17_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__39209\,
            in1 => \N__39631\,
            in2 => \N__34614\,
            in3 => \N__37822\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i19_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__37269\,
            in1 => \N__39675\,
            in2 => \N__29757\,
            in3 => \N__37824\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7_4_lut_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28044\,
            in1 => \N__28032\,
            in2 => \N__28021\,
            in3 => \N__28179\,
            lcout => OPEN,
            ltout => \ADC_VDC.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i11_3_lut_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28168\,
            in2 => \N__28159\,
            in3 => \N__28156\,
            lcout => \ADC_VDC.adc_state_3_N_1316_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19130_2_lut_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32849\,
            in2 => \_gnd_net_\,
            in3 => \N__32495\,
            lcout => \ADC_VDC.n22055\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i2_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32496\,
            in1 => \N__33273\,
            in2 => \_gnd_net_\,
            in3 => \N__33576\,
            lcout => adc_state_2_adj_1550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42753\,
            ce => \N__28141\,
            sr => \N__28108\
        );

    \ADC_VDC.i1_4_lut_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__28147\,
            in1 => \N__33575\,
            in2 => \N__33348\,
            in3 => \N__30517\,
            lcout => \ADC_VDC.n21871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i3_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011110000000"
        )
    port map (
            in0 => \N__33532\,
            in1 => \N__32485\,
            in2 => \N__33368\,
            in3 => \N__32599\,
            lcout => adc_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42717\,
            ce => \N__28132\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i14825_3_lut_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__32833\,
            in1 => \N__32450\,
            in2 => \_gnd_net_\,
            in3 => \N__33531\,
            lcout => OPEN,
            ltout => \ADC_VDC.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_15_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111010"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__28121\,
            in2 => \N__28126\,
            in3 => \N__32597\,
            lcout => \ADC_VDC.n44_adj_1487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i20180_3_lut_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__28122\,
            in2 => \_gnd_net_\,
            in3 => \N__32598\,
            lcout => \ADC_VDC.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100110010"
        )
    port map (
            in0 => \N__33314\,
            in1 => \N__33550\,
            in2 => \N__32848\,
            in3 => \N__32700\,
            lcout => \ADC_VDC.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42696\,
            ce => \N__30841\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33393\,
            in1 => \N__31082\,
            in2 => \N__33741\,
            in3 => \N__28438\,
            lcout => buf_adcdata_vdc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__28277\,
            in1 => \N__28426\,
            in2 => \N__28402\,
            in3 => \N__32701\,
            lcout => cmd_rdadctmp_9_adj_1565,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i11_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__31060\,
            in1 => \N__33354\,
            in2 => \N__28258\,
            in3 => \N__41241\,
            lcout => buf_adcdata_vdc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_adj_12_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001010000000"
        )
    port map (
            in0 => \N__32490\,
            in1 => \N__33551\,
            in2 => \N__33403\,
            in3 => \N__32688\,
            lcout => \ADC_VDC.n14120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31061\,
            in1 => \N__33355\,
            in2 => \N__35214\,
            in3 => \N__28243\,
            lcout => buf_adcdata_vdc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__33353\,
            in1 => \N__31063\,
            in2 => \N__28231\,
            in3 => \N__28206\,
            lcout => buf_adcdata_vdc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i16_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33352\,
            in1 => \N__31062\,
            in2 => \N__43536\,
            in3 => \N__28195\,
            lcout => buf_adcdata_vdc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i7_12609_12610_set_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36553\,
            in1 => \_gnd_net_\,
            in2 => \N__36187\,
            in3 => \N__31251\,
            lcout => \comm_spi.n15337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53691\,
            ce => 'H',
            sr => \N__41903\
        );

    \mux_126_Mux_5_i111_3_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36919\,
            in1 => \N__36940\,
            in2 => \_gnd_net_\,
            in3 => \N__59326\,
            lcout => n111_adj_1732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_5_i16_3_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59325\,
            in1 => \N__28723\,
            in2 => \_gnd_net_\,
            in3 => \N__32372\,
            lcout => n16_adj_1728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_6_i16_3_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59324\,
            in1 => \N__31323\,
            in2 => \_gnd_net_\,
            in3 => \N__31839\,
            lcout => n16_adj_1721,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_6_i19_3_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28696\,
            in1 => \N__28671\,
            in2 => \_gnd_net_\,
            in3 => \N__59323\,
            lcout => n19_adj_1722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i13037_2_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32696\,
            in2 => \_gnd_net_\,
            in3 => \N__28589\,
            lcout => \ADC_VDC.n15721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i5_12636_12637_reset_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28879\,
            in1 => \N__31456\,
            in2 => \_gnd_net_\,
            in3 => \N__33771\,
            lcout => \comm_spi.n15365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53690\,
            ce => 'H',
            sr => \N__35236\
        );

    \ADC_VDC.i1_3_lut_4_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110000000"
        )
    port map (
            in0 => \N__32509\,
            in1 => \N__33574\,
            in2 => \N__33439\,
            in3 => \N__32729\,
            lcout => \ADC_VDC.n14092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__28467\,
            in1 => \N__32508\,
            in2 => \_gnd_net_\,
            in3 => \N__30535\,
            lcout => OPEN,
            ltout => \ADC_VDC.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i34_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__33410\,
            in1 => \N__28483\,
            in2 => \N__28477\,
            in3 => \N__32730\,
            lcout => cmd_rdadcbuf_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42759\,
            ce => \N__28450\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_17_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__32507\,
            in1 => \N__33573\,
            in2 => \N__33438\,
            in3 => \N__32728\,
            lcout => n12352,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__36294\,
            in1 => \_gnd_net_\,
            in2 => \N__57147\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_857\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20238_4_lut_3_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28875\,
            in1 => \N__36295\,
            in2 => \_gnd_net_\,
            in3 => \N__57135\,
            lcout => \comm_spi.n24028\,
            ltout => \comm_spi.n24028_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i5_12636_12637_set_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__31452\,
            in1 => \_gnd_net_\,
            in2 => \N__28864\,
            in3 => \N__33772\,
            lcout => \comm_spi.n15364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53699\,
            ce => 'H',
            sr => \N__36157\
        );

    \comm_spi.i20243_4_lut_3_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36590\,
            in1 => \N__45657\,
            in2 => \_gnd_net_\,
            in3 => \N__57136\,
            lcout => \comm_spi.n24025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__57131\,
            in1 => \N__40657\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_854\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i20_3_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28861\,
            in1 => \N__28901\,
            in2 => \_gnd_net_\,
            in3 => \N__59327\,
            lcout => n20_adj_1781,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i20_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35958\,
            in1 => \N__28769\,
            in2 => \N__28825\,
            in3 => \N__33972\,
            lcout => cmd_rdadctmp_20_adj_1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23306_bdd_4_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__45601\,
            in1 => \N__43444\,
            in2 => \N__37462\,
            in3 => \N__60047\,
            lcout => n23309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19237_3_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28750\,
            in1 => \N__28940\,
            in2 => \_gnd_net_\,
            in3 => \N__59371\,
            lcout => OPEN,
            ltout => \n22164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20513_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__31462\,
            in1 => \N__60045\,
            in2 => \N__29071\,
            in3 => \N__60640\,
            lcout => n23468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i16_3_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29068\,
            in1 => \N__32235\,
            in2 => \_gnd_net_\,
            in3 => \N__59372\,
            lcout => OPEN,
            ltout => \n16_adj_1763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23366_bdd_4_lut_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__31630\,
            in1 => \N__29047\,
            in2 => \N__29035\,
            in3 => \N__60046\,
            lcout => n23369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_5_i127_3_lut_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36918\,
            in1 => \N__29026\,
            in2 => \_gnd_net_\,
            in3 => \N__61395\,
            lcout => \comm_buf_2_7_N_575_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i6_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__48808\,
            in1 => \N__57861\,
            in2 => \N__28994\,
            in3 => \N__40562\,
            lcout => \buf_cfgRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47452\,
            in1 => \N__48809\,
            in2 => \_gnd_net_\,
            in3 => \N__28941\,
            lcout => \buf_cfgRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i4_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48807\,
            in1 => \N__47373\,
            in2 => \_gnd_net_\,
            in3 => \N__28900\,
            lcout => \buf_cfgRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i12_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47374\,
            in1 => \N__50722\,
            in2 => \_gnd_net_\,
            in3 => \N__32282\,
            lcout => buf_dds0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i5_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__50723\,
            in1 => \N__56569\,
            in2 => \N__32376\,
            in3 => \N__57862\,
            lcout => buf_dds0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i19_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__57860\,
            in1 => \N__31431\,
            in2 => \N__62100\,
            in3 => \N__45421\,
            lcout => comm_test_buf_24_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i10_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39421\,
            in1 => \N__39732\,
            in2 => \N__29764\,
            in3 => \N__42056\,
            lcout => buf_adcdata_iac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i11_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__29732\,
            in1 => \N__55401\,
            in2 => \N__62101\,
            in3 => \N__49559\,
            lcout => buf_dds1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_count_i0_i0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29630\,
            in2 => \N__49437\,
            in3 => \_gnd_net_\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => n20613,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29522\,
            in2 => \_gnd_net_\,
            in3 => \N__29500\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n20613,
            carryout => n20614,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29414\,
            in2 => \_gnd_net_\,
            in3 => \N__29392\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n20614,
            carryout => n20615,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29309\,
            in2 => \_gnd_net_\,
            in3 => \N__29287\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n20615,
            carryout => n20616,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29198\,
            in2 => \_gnd_net_\,
            in3 => \N__29179\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n20616,
            carryout => n20617,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29096\,
            in2 => \_gnd_net_\,
            in3 => \N__29074\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n20617,
            carryout => n20618,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i6_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30161\,
            in2 => \_gnd_net_\,
            in3 => \N__30142\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n20618,
            carryout => n20619,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30053\,
            in2 => \_gnd_net_\,
            in3 => \N__30034\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n20619,
            carryout => n20620,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__50013\,
            sr => \N__49956\
        );

    \data_count_i0_i8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29951\,
            in2 => \_gnd_net_\,
            in3 => \N__29929\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => n20621,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__50019\,
            sr => \N__49957\
        );

    \data_count_i0_i9_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29846\,
            in2 => \_gnd_net_\,
            in3 => \N__29926\,
            lcout => data_count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__50019\,
            sr => \N__49957\
        );

    \i1_2_lut_4_lut_adj_270_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__55635\,
            in1 => \N__30560\,
            in2 => \N__38775\,
            in3 => \N__50887\,
            lcout => OPEN,
            ltout => \n24_adj_1598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__40940\,
            in1 => \N__29824\,
            in2 => \N__29815\,
            in3 => \N__43618\,
            lcout => \IAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61933\,
            ce => \N__36799\,
            sr => \N__37141\
        );

    \i1_2_lut_4_lut_adj_271_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__55636\,
            in1 => \N__29789\,
            in2 => \N__38776\,
            in3 => \N__50888\,
            lcout => OPEN,
            ltout => \n24_adj_1506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__62093\,
            in1 => \N__29770\,
            in2 => \N__29812\,
            in3 => \N__43423\,
            lcout => \IAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61933\,
            ce => \N__36799\,
            sr => \N__37141\
        );

    \i1_4_lut_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__59431\,
            in1 => \N__49322\,
            in2 => \N__46123\,
            in3 => \N__37394\,
            lcout => n11982,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_276_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__55634\,
            in1 => \N__38657\,
            in2 => \N__38774\,
            in3 => \N__50886\,
            lcout => n24_adj_1503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i16_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39377\,
            in1 => \N__39767\,
            in2 => \N__34385\,
            in3 => \N__30510\,
            lcout => buf_adcdata_iac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i6_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39766\,
            in1 => \N__32160\,
            in2 => \N__30490\,
            in3 => \N__37794\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23468_bdd_4_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__30469\,
            in1 => \N__30541\,
            in2 => \N__30619\,
            in3 => \N__60095\,
            lcout => n23471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i17_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39764\,
            in1 => \N__39378\,
            in2 => \N__30267\,
            in3 => \N__30456\,
            lcout => buf_adcdata_iac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_264_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31911\,
            in2 => \_gnd_net_\,
            in3 => \N__32147\,
            lcout => n13_adj_1591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.DTRIG_39_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101000"
        )
    port map (
            in0 => \N__30435\,
            in1 => \N__32148\,
            in2 => \N__30373\,
            in3 => \N__39768\,
            lcout => acadc_dtrig_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i28_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39765\,
            in1 => \N__37187\,
            in2 => \N__30304\,
            in3 => \N__37793\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20567_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__37047\,
            in1 => \N__60620\,
            in2 => \N__30263\,
            in3 => \N__59428\,
            lcout => n23534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i10_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31854\,
            in1 => \_gnd_net_\,
            in2 => \N__47453\,
            in3 => \N__50770\,
            lcout => buf_dds0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61967\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i15_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50771\,
            in1 => \N__57876\,
            in2 => \N__46663\,
            in3 => \N__32195\,
            lcout => buf_dds0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61967\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19233_3_lut_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30643\,
            in1 => \N__31853\,
            in2 => \_gnd_net_\,
            in3 => \N__59430\,
            lcout => n22160,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19234_3_lut_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59429\,
            in1 => \N__30599\,
            in2 => \_gnd_net_\,
            in3 => \N__30564\,
            lcout => n22161,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_9_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33249\,
            in2 => \_gnd_net_\,
            in3 => \N__32590\,
            lcout => \ADC_VDC.n21991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32591\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33266\,
            lcout => \ADC_VDC.n21707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_3__I_0_56_Mux_1_i10_3_lut_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100110"
        )
    port map (
            in0 => \N__32484\,
            in1 => \N__33581\,
            in2 => \_gnd_net_\,
            in3 => \N__30531\,
            lcout => \ADC_VDC.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i20026_4_lut_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__33086\,
            in1 => \N__30685\,
            in2 => \N__32641\,
            in3 => \N__32881\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i35_4_lut_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001010101"
        )
    port map (
            in0 => \N__32853\,
            in1 => \N__33151\,
            in2 => \N__30520\,
            in3 => \N__32457\,
            lcout => \ADC_VDC.n17\,
            ltout => \ADC_VDC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i33_3_lut_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32852\,
            in2 => \N__30715\,
            in3 => \N__33549\,
            lcout => OPEN,
            ltout => \ADC_VDC.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_14_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__30712\,
            in1 => \N__33318\,
            in2 => \N__30703\,
            in3 => \N__32595\,
            lcout => \ADC_VDC.n21869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i1_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__30700\,
            in1 => \N__33319\,
            in2 => \N__30661\,
            in3 => \N__32596\,
            lcout => adc_state_1_adj_1551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42698\,
            ce => \N__30694\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_6_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100000"
        )
    port map (
            in0 => \N__33534\,
            in1 => \N__32472\,
            in2 => \N__33429\,
            in3 => \N__32605\,
            lcout => \ADC_VDC.n13957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_13_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33115\,
            in2 => \_gnd_net_\,
            in3 => \N__30819\,
            lcout => \ADC_VDC.n11923\,
            ltout => \ADC_VDC.n11923_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_11_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30832\,
            in1 => \N__33146\,
            in2 => \N__30679\,
            in3 => \N__33008\,
            lcout => \ADC_VDC.n20869\,
            ltout => \ADC_VDC.n20869_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i5307_4_lut_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101101001100"
        )
    port map (
            in0 => \N__32470\,
            in1 => \N__33533\,
            in2 => \N__30676\,
            in3 => \N__32850\,
            lcout => \ADC_VDC.n8031\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.n23528_bdd_4_lut_4_lut_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100001100"
        )
    port map (
            in0 => \N__33536\,
            in1 => \N__30808\,
            in2 => \N__33430\,
            in3 => \N__33157\,
            lcout => \ADC_VDC.n23531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19149_2_lut_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33535\,
            in2 => \_gnd_net_\,
            in3 => \N__30649\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_16_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__30862\,
            in1 => \N__32471\,
            in2 => \N__30850\,
            in3 => \N__30847\,
            lcout => \ADC_VDC.n39_adj_1488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_10_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33066\,
            in2 => \_gnd_net_\,
            in3 => \N__33039\,
            lcout => \ADC_VDC.n6_adj_1485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__32961\,
            in1 => \N__32976\,
            in2 => \_gnd_net_\,
            in3 => \N__32943\,
            lcout => \ADC_VDC.n21859\,
            ltout => \ADC_VDC.n21859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_3_lut_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33116\,
            in2 => \N__30826\,
            in3 => \N__33144\,
            lcout => \ADC_VDC.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i20014_4_lut_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__33145\,
            in1 => \N__33117\,
            in2 => \N__33088\,
            in3 => \N__33040\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i20101_4_lut_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__33548\,
            in1 => \N__33007\,
            in2 => \N__30823\,
            in3 => \N__30820\,
            lcout => \ADC_VDC.n22625\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__33041\,
            in1 => \N__33006\,
            in2 => \N__33087\,
            in3 => \N__30802\,
            lcout => \ADC_VDC.n11183\,
            ltout => \ADC_VDC.n11183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i23_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__30753\,
            in1 => \N__30796\,
            in2 => \N__30763\,
            in3 => \N__32494\,
            lcout => \ADC_VDC.cmd_rdadctmp_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42697\,
            ce => \N__30739\,
            sr => \N__30724\
        );

    \comm_spi.imiso_83_12612_12613_reset_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38181\,
            in1 => \N__38436\,
            in2 => \_gnd_net_\,
            in3 => \N__41986\,
            lcout => \comm_spi.n15341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12612_12613_resetC_net\,
            ce => 'H',
            sr => \N__40629\
        );

    \comm_spi.data_tx_i7_12609_12610_reset_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36183\,
            in1 => \N__31252\,
            in2 => \_gnd_net_\,
            in3 => \N__36552\,
            lcout => \comm_spi.n15338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53666\,
            ce => 'H',
            sr => \N__40630\
        );

    \comm_cmd_1__bdd_4_lut_20473_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__59328\,
            in1 => \N__31234\,
            in2 => \N__31114\,
            in3 => \N__60544\,
            lcout => OPEN,
            ltout => \n23384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23384_bdd_4_lut_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__31197\,
            in1 => \N__31170\,
            in2 => \N__31135\,
            in3 => \N__59330\,
            lcout => n23387,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i21_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31033\,
            in1 => \N__33387\,
            in2 => \N__31113\,
            in3 => \N__31132\,
            lcout => buf_adcdata_vdc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i13_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__33385\,
            in1 => \N__31099\,
            in2 => \N__31073\,
            in3 => \N__38061\,
            lcout => buf_adcdata_vdc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31032\,
            in1 => \N__33386\,
            in2 => \N__37899\,
            in3 => \N__30964\,
            lcout => buf_adcdata_vdc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_4_i19_3_lut_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30946\,
            in1 => \N__30918\,
            in2 => \_gnd_net_\,
            in3 => \N__59329\,
            lcout => OPEN,
            ltout => \n19_adj_1734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20498_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__30889\,
            in1 => \N__60036\,
            in2 => \N__30865\,
            in3 => \N__60545\,
            lcout => n23438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_124_Mux_1_i30_4_lut_4_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111011001"
        )
    port map (
            in0 => \N__60546\,
            in1 => \N__61032\,
            in2 => \N__60090\,
            in3 => \N__59331\,
            lcout => n30_adj_1805,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i8_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35999\,
            in1 => \N__36113\,
            in2 => \N__31393\,
            in3 => \N__34002\,
            lcout => cmd_rdadctmp_8_adj_1540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i7_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33990\,
            in1 => \N__31389\,
            in2 => \N__31381\,
            in3 => \N__36001\,
            lcout => cmd_rdadctmp_7_adj_1541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i6_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__35998\,
            in1 => \N__33991\,
            in2 => \N__31369\,
            in3 => \N__31377\,
            lcout => cmd_rdadctmp_6_adj_1542,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i5_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33989\,
            in1 => \N__31365\,
            in2 => \N__31339\,
            in3 => \N__36000\,
            lcout => cmd_rdadctmp_5_adj_1543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35997\,
            in1 => \N__31335\,
            in2 => \N__34006\,
            in3 => \N__31356\,
            lcout => cmd_rdadctmp_4_adj_1544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i6_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__31322\,
            in1 => \N__55399\,
            in2 => \N__49243\,
            in3 => \N__49503\,
            lcout => buf_dds1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i9_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__35421\,
            in1 => \N__38128\,
            in2 => \N__39807\,
            in3 => \N__37840\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_0_i30_3_lut_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31300\,
            in1 => \N__60989\,
            in2 => \_gnd_net_\,
            in3 => \N__37855\,
            lcout => n30_adj_1588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i13_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35616\,
            in1 => \N__35962\,
            in2 => \N__31282\,
            in3 => \N__38036\,
            lcout => buf_adcdata_vac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_7_i127_3_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__61396\,
            in1 => \N__38352\,
            in2 => \_gnd_net_\,
            in3 => \N__31567\,
            lcout => \comm_buf_2_7_N_575_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i17_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35617\,
            in1 => \N__35963\,
            in2 => \N__31555\,
            in3 => \N__48602\,
            lcout => buf_adcdata_vac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i20_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__57863\,
            in1 => \N__31417\,
            in2 => \N__44707\,
            in3 => \N__45414\,
            lcout => comm_test_buf_24_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19236_3_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31516\,
            in1 => \N__31485\,
            in2 => \_gnd_net_\,
            in3 => \N__59020\,
            lcout => n22163,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_12632_12633_set_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36238\,
            in1 => \N__34045\,
            in2 => \_gnd_net_\,
            in3 => \N__51052\,
            lcout => \comm_spi.n15360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53710\,
            ce => 'H',
            sr => \N__31441\
        );

    \mux_125_Mux_3_i111_3_lut_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31432\,
            in1 => \N__34257\,
            in2 => \_gnd_net_\,
            in3 => \N__59261\,
            lcout => n111_adj_1794,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_3_i111_3_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__59262\,
            in1 => \N__34178\,
            in2 => \_gnd_net_\,
            in3 => \N__34258\,
            lcout => n111_adj_1744,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i111_3_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59263\,
            in1 => \N__31416\,
            in2 => \_gnd_net_\,
            in3 => \N__34245\,
            lcout => n111_adj_1785,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_4_i111_3_lut_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__59264\,
            in1 => \N__34091\,
            in2 => \_gnd_net_\,
            in3 => \N__34246\,
            lcout => n111_adj_1737,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_289_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__50893\,
            in1 => \N__31644\,
            in2 => \N__55651\,
            in3 => \N__38757\,
            lcout => OPEN,
            ltout => \n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__31573\,
            in1 => \N__40561\,
            in2 => \N__31693\,
            in3 => \N__43611\,
            lcout => \VAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61872\,
            ce => \N__36798\,
            sr => \N__37126\
        );

    \mux_125_Mux_6_i17_3_lut_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31683\,
            in1 => \N__31643\,
            in2 => \_gnd_net_\,
            in3 => \N__59265\,
            lcout => n17_adj_1764,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_64_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__59267\,
            in1 => \N__55822\,
            in2 => \N__40429\,
            in3 => \N__37405\,
            lcout => OPEN,
            ltout => \n11981_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__46621\,
            in1 => \N__31579\,
            in2 => \N__31621\,
            in3 => \N__43422\,
            lcout => \VAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61872\,
            ce => \N__36798\,
            sr => \N__37126\
        );

    \i1_2_lut_4_lut_adj_292_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__55626\,
            in1 => \N__50892\,
            in2 => \N__38772\,
            in3 => \N__31595\,
            lcout => n24_adj_1576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_57_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__37404\,
            in1 => \N__49214\,
            in2 => \N__36346\,
            in3 => \N__59266\,
            lcout => n11986,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10511_3_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40425\,
            in1 => \N__46620\,
            in2 => \_gnd_net_\,
            in3 => \N__46202\,
            lcout => n13237,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20548_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__60041\,
            in1 => \N__60587\,
            in2 => \N__50221\,
            in3 => \N__31723\,
            lcout => OPEN,
            ltout => \n23510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23510_bdd_4_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__41482\,
            in1 => \N__44365\,
            in2 => \N__31741\,
            in3 => \N__60042\,
            lcout => OPEN,
            ltout => \n23513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1663271_i1_3_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31738\,
            in2 => \N__31729\,
            in3 => \N__61055\,
            lcout => OPEN,
            ltout => \n30_adj_1759_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_7_i127_3_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31708\,
            in2 => \N__31726\,
            in3 => \N__61397\,
            lcout => \comm_buf_0_7_N_543_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_7_i26_3_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47293\,
            in1 => \N__59268\,
            in2 => \_gnd_net_\,
            in3 => \N__31716\,
            lcout => n26_adj_1758,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_302_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__31717\,
            in1 => \N__39173\,
            in2 => \N__34705\,
            in3 => \N__31699\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_end_302C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_7_i112_3_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38351\,
            in1 => \N__36880\,
            in2 => \_gnd_net_\,
            in3 => \N__60588\,
            lcout => n112_adj_1762,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110000101100"
        )
    port map (
            in0 => \N__45787\,
            in1 => \N__34782\,
            in2 => \N__34699\,
            in3 => \N__49435\,
            lcout => n17_adj_1742,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_272_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__45781\,
            in1 => \N__31762\,
            in2 => \N__34796\,
            in3 => \N__34274\,
            lcout => OPEN,
            ltout => \n21946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20133_3_lut_4_lut_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__34783\,
            in1 => \N__45782\,
            in2 => \N__31702\,
            in3 => \N__34685\,
            lcout => n21880,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i34_3_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49436\,
            in1 => \N__34784\,
            in2 => \_gnd_net_\,
            in3 => \N__41370\,
            lcout => OPEN,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__45790\,
            in1 => \N__34686\,
            in2 => \N__31810\,
            in3 => \N__31807\,
            lcout => eis_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i2C_net\,
            ce => \N__34423\,
            sr => \N__39178\
        );

    \i19812_2_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34275\,
            lcout => n22395,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20187_2_lut_3_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__45788\,
            in1 => \_gnd_net_\,
            in2 => \N__34698\,
            in3 => \N__39171\,
            lcout => n22120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20166_3_lut_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__31747\,
            in1 => \N__34678\,
            in2 => \_gnd_net_\,
            in3 => \N__45789\,
            lcout => n12369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i21_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39772\,
            in1 => \N__39398\,
            in2 => \N__32122\,
            in3 => \N__38606\,
            lcout => buf_adcdata_iac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i3_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110000"
        )
    port map (
            in0 => \N__48943\,
            in1 => \N__63778\,
            in2 => \N__55400\,
            in3 => \N__36860\,
            lcout => buf_dds1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i30_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39773\,
            in1 => \N__31778\,
            in2 => \N__32121\,
            in3 => \N__37836\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19796_2_lut_3_lut_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32146\,
            in2 => \N__31918\,
            in3 => \N__34672\,
            lcout => n22312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_265_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__43843\,
            in1 => \N__31761\,
            in2 => \N__34791\,
            in3 => \N__38872\,
            lcout => n11_adj_1592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i7_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__39774\,
            in1 => \N__32161\,
            in2 => \N__38160\,
            in3 => \N__37837\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_206_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__34671\,
            in1 => \N__31914\,
            in2 => \N__32149\,
            in3 => \_gnd_net_\,
            lcout => n17633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_adj_49_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31912\,
            in2 => \_gnd_net_\,
            in3 => \N__32142\,
            lcout => \iac_raw_buf_N_823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i7_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47521\,
            in1 => \N__50754\,
            in2 => \_gnd_net_\,
            in3 => \N__32312\,
            lcout => buf_dds0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i29_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__37188\,
            in2 => \N__39808\,
            in3 => \N__37795\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.DTRIG_39_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101000"
        )
    port map (
            in0 => \N__31913\,
            in1 => \N__32101\,
            in2 => \N__32011\,
            in3 => \N__36002\,
            lcout => acadc_dtrig_v,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23534_bdd_4_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__31890\,
            in1 => \N__31861\,
            in2 => \N__50644\,
            in3 => \N__60564\,
            lcout => n22177,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i10_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__50549\,
            in1 => \N__31855\,
            in2 => \N__32332\,
            in3 => \N__50415\,
            lcout => \SIG_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i6_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50552\,
            in1 => \N__50414\,
            in2 => \N__32341\,
            in3 => \N__31840\,
            lcout => \SIG_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50550\,
            in1 => \N__50413\,
            in2 => \N__37438\,
            in3 => \N__47269\,
            lcout => \SIG_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__50411\,
            in1 => \N__50551\,
            in2 => \N__32380\,
            in3 => \N__32347\,
            lcout => \SIG_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i9_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__50640\,
            in1 => \N__50554\,
            in2 => \N__32170\,
            in3 => \N__50416\,
            lcout => \SIG_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50412\,
            in1 => \N__50553\,
            in2 => \N__32323\,
            in3 => \N__32313\,
            lcout => \SIG_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61950\,
            ce => \N__42208\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i12_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__50544\,
            in1 => \N__50407\,
            in2 => \N__32293\,
            in3 => \N__32887\,
            lcout => \SIG_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61968\,
            ce => \N__42206\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i13_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50545\,
            in1 => \N__50408\,
            in2 => \N__32260\,
            in3 => \N__55549\,
            lcout => \SIG_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61968\,
            ce => \N__42206\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i14_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50546\,
            in1 => \N__50409\,
            in2 => \N__32251\,
            in3 => \N__32242\,
            lcout => \SIG_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61968\,
            ce => \N__42206\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i15_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50547\,
            in1 => \N__50410\,
            in2 => \N__32212\,
            in3 => \N__32196\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61968\,
            ce => \N__42206\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i8_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__50406\,
            in1 => \N__50548\,
            in2 => \N__40236\,
            in3 => \N__32176\,
            lcout => \SIG_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61968\,
            ce => \N__42206\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i11_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50543\,
            in1 => \N__50403\,
            in2 => \N__32923\,
            in3 => \N__32911\,
            lcout => \SIG_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61982\,
            ce => \N__42207\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19141_2_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32854\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33577\,
            lcout => \ADC_VDC.n22067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19137_2_lut_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \_gnd_net_\,
            in3 => \N__33043\,
            lcout => \ADC_VDC.n22063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35096\,
            in1 => \N__35061\,
            in2 => \_gnd_net_\,
            in3 => \N__35080\,
            lcout => \RTD.n20050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_7_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33579\,
            in2 => \_gnd_net_\,
            in3 => \N__32851\,
            lcout => OPEN,
            ltout => \ADC_VDC.n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i14816_4_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010000"
        )
    port map (
            in0 => \N__32702\,
            in1 => \N__32749\,
            in2 => \N__32752\,
            in3 => \N__33379\,
            lcout => \ADC_VDC.n17542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_8_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33578\,
            in2 => \_gnd_net_\,
            in3 => \N__32459\,
            lcout => \ADC_VDC.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i24_4_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001110010"
        )
    port map (
            in0 => \N__33378\,
            in1 => \N__32460\,
            in2 => \N__32743\,
            in3 => \N__32703\,
            lcout => \ADC_VDC.n17565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001101010"
        )
    port map (
            in0 => \N__32458\,
            in1 => \N__33580\,
            in2 => \N__33431\,
            in3 => \N__33163\,
            lcout => \ADC_VDC.n23528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.bit_cnt_3791__i0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33150\,
            in2 => \_gnd_net_\,
            in3 => \N__33121\,
            lcout => \ADC_VDC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \ADC_VDC.n20812\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33118\,
            in2 => \_gnd_net_\,
            in3 => \N__33091\,
            lcout => \ADC_VDC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20812\,
            carryout => \ADC_VDC.n20813\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33076\,
            in2 => \_gnd_net_\,
            in3 => \N__33046\,
            lcout => \ADC_VDC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20813\,
            carryout => \ADC_VDC.n20814\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33042\,
            in2 => \_gnd_net_\,
            in3 => \N__33013\,
            lcout => \ADC_VDC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20814\,
            carryout => \ADC_VDC.n20815\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33009\,
            in2 => \_gnd_net_\,
            in3 => \N__32980\,
            lcout => \ADC_VDC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20815\,
            carryout => \ADC_VDC.n20816\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32977\,
            in2 => \_gnd_net_\,
            in3 => \N__32965\,
            lcout => \ADC_VDC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20816\,
            carryout => \ADC_VDC.n20817\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32962\,
            in2 => \_gnd_net_\,
            in3 => \N__32950\,
            lcout => \ADC_VDC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n20817\,
            carryout => \ADC_VDC.n20818\,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \ADC_VDC.bit_cnt_3791__i7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32944\,
            in2 => \_gnd_net_\,
            in3 => \N__32947\,
            lcout => \ADC_VDC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42690\,
            ce => \N__32932\,
            sr => \N__33781\
        );

    \comm_spi.data_tx_i4_12632_12633_reset_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34035\,
            in1 => \N__36231\,
            in2 => \_gnd_net_\,
            in3 => \N__51045\,
            lcout => \comm_spi.n15361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53602\,
            ce => 'H',
            sr => \N__36274\
        );

    \mux_127_Mux_3_i19_3_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33748\,
            in1 => \N__33644\,
            in2 => \_gnd_net_\,
            in3 => \N__59398\,
            lcout => OPEN,
            ltout => \n19_adj_1703_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_3_i22_3_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33689\,
            in2 => \N__33724\,
            in3 => \N__60008\,
            lcout => OPEN,
            ltout => \n22_adj_1704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_3_i30_3_lut_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33721\,
            in2 => \N__33703\,
            in3 => \N__61013\,
            lcout => n30_adj_1705,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35625\,
            in1 => \N__35927\,
            in2 => \N__33805\,
            in3 => \N__33606\,
            lcout => buf_adcdata_vac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__33690\,
            in1 => \N__39404\,
            in2 => \N__35388\,
            in3 => \N__39817\,
            lcout => buf_adcdata_iac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__33645\,
            in1 => \N__35928\,
            in2 => \N__35629\,
            in3 => \N__33676\,
            lcout => buf_adcdata_vac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_4_lut_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__54609\,
            in1 => \N__64079\,
            in2 => \N__54424\,
            in3 => \N__63076\,
            lcout => n8_adj_1755,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_1_i19_3_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33631\,
            in1 => \N__33602\,
            in2 => \_gnd_net_\,
            in3 => \N__59250\,
            lcout => OPEN,
            ltout => \n19_adj_1710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_1_i22_3_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36086\,
            in2 => \N__34066\,
            in3 => \N__60040\,
            lcout => OPEN,
            ltout => \n22_adj_1711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_1_i30_3_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34063\,
            in2 => \N__34051\,
            in3 => \N__61056\,
            lcout => OPEN,
            ltout => \n30_adj_1712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_1_i127_3_lut_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41867\,
            in2 => \N__34048\,
            in3 => \N__61398\,
            lcout => \comm_buf_2_7_N_575_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20233_4_lut_3_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34023\,
            in1 => \N__57177\,
            in2 => \_gnd_net_\,
            in3 => \N__46078\,
            lcout => \comm_spi.n24031\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_3_i127_3_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34186\,
            in1 => \N__34012\,
            in2 => \_gnd_net_\,
            in3 => \N__61399\,
            lcout => \comm_buf_2_7_N_575_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i9_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35990\,
            in1 => \N__33797\,
            in2 => \N__36126\,
            in3 => \N__33993\,
            lcout => cmd_rdadctmp_9_adj_1539,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i10_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33992\,
            in1 => \N__36029\,
            in2 => \N__33804\,
            in3 => \N__35991\,
            lcout => cmd_rdadctmp_10_adj_1538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_6_i2_3_lut_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36342\,
            in1 => \N__40753\,
            in2 => \_gnd_net_\,
            in3 => \N__54422\,
            lcout => OPEN,
            ltout => \n2_adj_1666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__54611\,
            in1 => \N__34123\,
            in2 => \N__33784\,
            in3 => \N__34204\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61840\,
            ce => \N__46426\,
            sr => \N__46348\
        );

    \i20030_2_lut_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37990\,
            in2 => \_gnd_net_\,
            in3 => \N__54420\,
            lcout => n22295,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_6_i4_3_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54421\,
            in1 => \N__43126\,
            in2 => \_gnd_net_\,
            in3 => \N__53800\,
            lcout => n4_adj_1667,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_6_i1_3_lut_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49239\,
            in1 => \N__40503\,
            in2 => \_gnd_net_\,
            in3 => \N__54423\,
            lcout => n1_adj_1665,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10505_3_lut_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36341\,
            in1 => \N__40517\,
            in2 => \_gnd_net_\,
            in3 => \N__46204\,
            lcout => n13231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57178\,
            in2 => \_gnd_net_\,
            in3 => \N__36200\,
            lcout => \comm_spi.data_tx_7__N_865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__52144\,
            in2 => \_gnd_net_\,
            in3 => \N__38278\,
            lcout => comm_test_buf_24_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52936\,
            in1 => \N__36697\,
            in2 => \_gnd_net_\,
            in3 => \N__40867\,
            lcout => comm_test_buf_24_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i4_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36695\,
            in1 => \_gnd_net_\,
            in2 => \N__56109\,
            in3 => \N__36301\,
            lcout => comm_test_buf_24_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i6_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49230\,
            in1 => \N__36699\,
            in2 => \_gnd_net_\,
            in3 => \N__34072\,
            lcout => comm_test_buf_24_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i7_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__55848\,
            in2 => \_gnd_net_\,
            in3 => \N__34237\,
            lcout => comm_test_buf_24_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__43198\,
            in1 => \_gnd_net_\,
            in2 => \N__49141\,
            in3 => \N__36700\,
            lcout => comm_test_buf_24_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36694\,
            in1 => \N__49326\,
            in2 => \_gnd_net_\,
            in3 => \N__46093\,
            lcout => comm_test_buf_24_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \comm_test_buf_24_i5_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__56587\,
            in1 => \N__36698\,
            in2 => \_gnd_net_\,
            in3 => \N__37969\,
            lcout => comm_test_buf_24_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61846\,
            ce => \N__41188\,
            sr => \N__34156\
        );

    \n23324_bdd_4_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__34136\,
            in1 => \N__34354\,
            in2 => \N__40240\,
            in3 => \N__60462\,
            lcout => n23327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20419_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__54610\,
            in1 => \N__34228\,
            in2 => \N__34216\,
            in3 => \N__51837\,
            lcout => n23294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_0_i127_3_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48986\,
            in1 => \N__34195\,
            in2 => \_gnd_net_\,
            in3 => \N__61400\,
            lcout => \comm_buf_2_7_N_575_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i112_3_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60461\,
            in1 => \N__34179\,
            in2 => \_gnd_net_\,
            in3 => \N__34162\,
            lcout => n112_adj_1795,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12822_2_lut_3_lut_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__64097\,
            in1 => \N__41187\,
            in2 => \_gnd_net_\,
            in3 => \N__62607\,
            lcout => n15545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i8_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__55430\,
            in1 => \N__43955\,
            in2 => \N__34143\,
            in3 => \N__49537\,
            lcout => buf_dds1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12815_2_lut_3_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__36777\,
            in1 => \N__62603\,
            in2 => \_gnd_net_\,
            in3 => \N__64096\,
            lcout => n15538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i8_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43939\,
            in1 => \N__49106\,
            in2 => \_gnd_net_\,
            in3 => \N__36671\,
            lcout => comm_test_buf_24_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i11_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36665\,
            in1 => \N__62086\,
            in2 => \_gnd_net_\,
            in3 => \N__49318\,
            lcout => comm_test_buf_24_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i13_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45335\,
            in1 => \N__56583\,
            in2 => \_gnd_net_\,
            in3 => \N__36669\,
            lcout => comm_test_buf_24_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i9_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__52138\,
            in1 => \_gnd_net_\,
            in2 => \N__44630\,
            in3 => \N__36692\,
            lcout => comm_test_buf_24_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i10_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52934\,
            in1 => \N__40935\,
            in2 => \_gnd_net_\,
            in3 => \N__36668\,
            lcout => comm_test_buf_24_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i12_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36666\,
            in1 => \N__44703\,
            in2 => \_gnd_net_\,
            in3 => \N__56110\,
            lcout => comm_test_buf_24_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i14_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49231\,
            in1 => \N__40539\,
            in2 => \_gnd_net_\,
            in3 => \N__36670\,
            lcout => comm_test_buf_24_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_test_buf_24_i15_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36667\,
            in1 => \_gnd_net_\,
            in2 => \N__46629\,
            in3 => \N__55823\,
            lcout => comm_test_buf_24_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61862\,
            ce => \N__44044\,
            sr => \N__41338\
        );

    \comm_cmd_0__bdd_4_lut_20562_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__34343\,
            in1 => \N__60589\,
            in2 => \N__43842\,
            in3 => \N__59113\,
            lcout => n23522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20409_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__59114\,
            in1 => \N__34386\,
            in2 => \N__37083\,
            in3 => \N__60627\,
            lcout => n23324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34344\,
            in1 => \N__48870\,
            in2 => \_gnd_net_\,
            in3 => \N__51361\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_256_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__49756\,
            in1 => \N__50065\,
            in2 => \N__34345\,
            in3 => \N__60689\,
            lcout => OPEN,
            ltout => \n19_adj_1727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44056\,
            in1 => \N__44128\,
            in2 => \N__34327\,
            in3 => \N__38452\,
            lcout => OPEN,
            ltout => \n29_adj_1770_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38867\,
            in2 => \N__34324\,
            in3 => \N__41464\,
            lcout => n16_adj_1683,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__60690\,
            in1 => \N__55276\,
            in2 => \_gnd_net_\,
            in3 => \N__51360\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_6_i111_3_lut_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__59115\,
            in1 => \_gnd_net_\,
            in2 => \N__34320\,
            in3 => \N__34293\,
            lcout => n111_adj_1726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14917_4_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__43835\,
            in1 => \N__34276\,
            in2 => \N__34695\,
            in3 => \N__41551\,
            lcout => OPEN,
            ltout => \n17642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000010001"
        )
    port map (
            in0 => \N__34774\,
            in1 => \N__34670\,
            in2 => \N__34261\,
            in3 => \N__34555\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__34419\,
            sr => \N__39172\
        );

    \eis_state_1__bdd_4_lut_4_lut_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101011101010"
        )
    port map (
            in0 => \N__45797\,
            in1 => \N__34561\,
            in2 => \N__34786\,
            in3 => \N__34548\,
            lcout => n23330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3823_3_lut_3_lut_4_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__45798\,
            in1 => \N__39132\,
            in2 => \N__34787\,
            in3 => \N__34549\,
            lcout => \iac_raw_buf_N_821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_4_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__34666\,
            in1 => \N__45783\,
            in2 => \N__34785\,
            in3 => \N__39131\,
            lcout => n12394,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__34429\,
            in1 => \N__45799\,
            in2 => \N__34795\,
            in3 => \N__41371\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__34419\,
            sr => \N__39172\
        );

    \buf_device_acadc_i2_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__37018\,
            in1 => \N__34804\,
            in2 => \N__44647\,
            in3 => \N__43617\,
            lcout => \IAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61901\,
            ce => \N__36790\,
            sr => \N__37134\
        );

    \buf_device_acadc_i6_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__43616\,
            in1 => \N__45326\,
            in2 => \N__34402\,
            in3 => \N__37012\,
            lcout => \VAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61901\,
            ce => \N__36790\,
            sr => \N__37134\
        );

    \i16467_2_lut_3_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__64109\,
            in1 => \N__52107\,
            in2 => \_gnd_net_\,
            in3 => \N__62604\,
            lcout => n14_adj_1613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16445_2_lut_3_lut_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__64111\,
            in1 => \N__56570\,
            in2 => \_gnd_net_\,
            in3 => \N__62605\,
            lcout => n14_adj_1661,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_77_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45325\,
            in1 => \N__62606\,
            in2 => \_gnd_net_\,
            in3 => \N__64110\,
            lcout => n14_adj_1660,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_335_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__52143\,
            in1 => \N__37382\,
            in2 => \N__59514\,
            in3 => \N__38311\,
            lcout => n11980,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i9_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63526\,
            in1 => \N__44515\,
            in2 => \N__57747\,
            in3 => \N__44497\,
            lcout => data_index_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20191_3_lut_4_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__45800\,
            in1 => \N__34696\,
            in2 => \N__34797\,
            in3 => \N__39130\,
            lcout => n12450,
            ltout => \n12450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20174_2_lut_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__34697\,
            in1 => \_gnd_net_\,
            in2 => \N__34618\,
            in3 => \_gnd_net_\,
            lcout => n15439,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i12_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39762\,
            in1 => \N__39370\,
            in2 => \N__37254\,
            in3 => \N__36977\,
            lcout => buf_adcdata_iac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i21_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57661\,
            in1 => \N__45327\,
            in2 => \N__36955\,
            in3 => \N__45426\,
            lcout => comm_test_buf_24_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i8_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39763\,
            in1 => \N__39371\,
            in2 => \N__34615\,
            in3 => \N__46946\,
            lcout => buf_adcdata_iac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49412\,
            in2 => \N__39982\,
            in3 => \_gnd_net_\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => n20637,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__35171\,
            sr => \N__34573\
        );

    \add_70_2_THRU_CRY_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64807\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n20637,
            carryout => \n20637_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_1_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__64852\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_0_THRU_CO\,
            carryout => \n20637_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_2_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64811\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_1_THRU_CO\,
            carryout => \n20637_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_3_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__64853\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_2_THRU_CO\,
            carryout => \n20637_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_4_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64815\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_3_THRU_CO\,
            carryout => \n20637_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_5_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__64854\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_4_THRU_CO\,
            carryout => \n20637_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_70_2_THRU_CRY_6_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64819\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n20637_THRU_CRY_5_THRU_CO\,
            carryout => \n20637_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44010\,
            in2 => \_gnd_net_\,
            in3 => \N__34813\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => n20638,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i2_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38961\,
            in2 => \_gnd_net_\,
            in3 => \N__34810\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n20638,
            carryout => n20639,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i3_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41526\,
            in2 => \_gnd_net_\,
            in3 => \N__34807\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n20639,
            carryout => n20640,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i4_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43986\,
            in2 => \_gnd_net_\,
            in3 => \N__34840\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n20640,
            carryout => n20641,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i5_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41157\,
            in2 => \_gnd_net_\,
            in3 => \N__34837\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n20641,
            carryout => n20642,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i6_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39957\,
            in2 => \_gnd_net_\,
            in3 => \N__34834\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n20642,
            carryout => n20643,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i7_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38979\,
            in2 => \_gnd_net_\,
            in3 => \N__34831\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n20643,
            carryout => n20644,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i8_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41601\,
            in2 => \_gnd_net_\,
            in3 => \N__34828\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n20644,
            carryout => n20645,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__35188\,
            sr => \N__35154\
        );

    \acadc_skipcnt_i0_i9_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37329\,
            in2 => \_gnd_net_\,
            in3 => \N__34825\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => n20646,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i10_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38925\,
            in2 => \_gnd_net_\,
            in3 => \N__34822\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n20646,
            carryout => n20647,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i11_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37299\,
            in2 => \_gnd_net_\,
            in3 => \N__34819\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n20647,
            carryout => n20648,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i12_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38943\,
            in2 => \_gnd_net_\,
            in3 => \N__34816\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n20648,
            carryout => n20649,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i13_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38835\,
            in2 => \_gnd_net_\,
            in3 => \N__35197\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n20649,
            carryout => n20650,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i14_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37314\,
            in2 => \_gnd_net_\,
            in3 => \N__35194\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n20650,
            carryout => n20651,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \acadc_skipcnt_i0_i15_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37347\,
            in2 => \_gnd_net_\,
            in3 => \N__35191\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__35187\,
            sr => \N__35155\
        );

    \clk_RTD_290_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__34885\,
            in1 => \N__36465\,
            in2 => \_gnd_net_\,
            in3 => \N__36439\,
            lcout => \clk_RTD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3789__i3_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__35065\,
            in1 => \N__35117\,
            in2 => \N__35101\,
            in3 => \N__35083\,
            lcout => \RTD.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34886\,
            ce => \N__34864\,
            sr => \N__34852\
        );

    \RTD.bit_cnt_3789__i2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__35082\,
            in1 => \N__35097\,
            in2 => \_gnd_net_\,
            in3 => \N__35064\,
            lcout => \RTD.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34886\,
            ce => \N__34864\,
            sr => \N__34852\
        );

    \RTD.bit_cnt_3789__i1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35081\,
            lcout => \RTD.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34886\,
            ce => \N__34864\,
            sr => \N__34852\
        );

    \RTD.bit_cnt_3789__i0_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35062\,
            lcout => \RTD.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34886\,
            ce => \N__34864\,
            sr => \N__34852\
        );

    \clk_cnt_3781_3782__i2_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36437\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36458\,
            lcout => clk_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \N__36415\
        );

    \clk_cnt_3781_3782__i1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36436\,
            lcout => clk_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \N__36415\
        );

    \comm_cmd_0__bdd_4_lut_20518_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__35344\,
            in1 => \N__60590\,
            in2 => \N__35311\,
            in3 => \N__59397\,
            lcout => n23432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_257_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__57740\,
            in1 => \N__51396\,
            in2 => \N__42781\,
            in3 => \N__63649\,
            lcout => n12610,
            ltout => \n12610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i5_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__45312\,
            in1 => \N__57741\,
            in2 => \N__35275\,
            in3 => \N__36500\,
            lcout => \AMPV_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_2_lut_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__57137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43277\,
            lcout => \comm_spi.data_tx_7__N_883\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12608_3_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41981\,
            in1 => \N__37492\,
            in2 => \_gnd_net_\,
            in3 => \N__41935\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_308_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__64065\,
            in1 => \N__63648\,
            in2 => \N__62677\,
            in3 => \N__63047\,
            lcout => n13117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45653\,
            in2 => \_gnd_net_\,
            in3 => \N__57109\,
            lcout => \comm_spi.data_tx_7__N_868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_2_i19_3_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35221\,
            in1 => \N__35447\,
            in2 => \_gnd_net_\,
            in3 => \N__59181\,
            lcout => OPEN,
            ltout => \n19_adj_1706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_2_i22_3_lut_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36056\,
            in2 => \N__36130\,
            in3 => \N__60007\,
            lcout => n22_adj_1707,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35623\,
            in1 => \N__35929\,
            in2 => \N__36127\,
            in3 => \N__37878\,
            lcout => buf_adcdata_vac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39419\,
            in1 => \N__39812\,
            in2 => \N__36093\,
            in3 => \N__35433\,
            lcout => buf_adcdata_iac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__36057\,
            in1 => \N__35409\,
            in2 => \N__39820\,
            in3 => \N__39420\,
            lcout => buf_adcdata_iac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__35448\,
            in1 => \N__36033\,
            in2 => \N__35989\,
            in3 => \N__35624\,
            lcout => buf_adcdata_vac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i10_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39811\,
            in1 => \N__35405\,
            in2 => \N__35434\,
            in3 => \N__37839\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i11_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37838\,
            in1 => \N__35378\,
            in2 => \N__35410\,
            in3 => \N__39816\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57172\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46071\,
            lcout => \comm_spi.data_tx_7__N_858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20228_4_lut_3_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51114\,
            in1 => \N__40855\,
            in2 => \_gnd_net_\,
            in3 => \N__57174\,
            lcout => \comm_spi.n24034\,
            ltout => \comm_spi.n24034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12628_12629_set_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51093\,
            in2 => \N__36241\,
            in3 => \N__51075\,
            lcout => \comm_spi.n15356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53627\,
            ce => 'H',
            sr => \N__36214\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40854\,
            in2 => \_gnd_net_\,
            in3 => \N__57173\,
            lcout => \comm_spi.data_tx_7__N_859\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57170\,
            lcout => \comm_spi.data_tx_7__N_855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20248_4_lut_3_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57175\,
            in1 => \N__36202\,
            in2 => \_gnd_net_\,
            in3 => \N__36168\,
            lcout => \comm_spi.n24013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45658\,
            in2 => \_gnd_net_\,
            in3 => \N__57171\,
            lcout => \comm_spi.data_tx_7__N_856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_4_i2_3_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36834\,
            in1 => \N__40699\,
            in2 => \_gnd_net_\,
            in3 => \N__54416\,
            lcout => OPEN,
            ltout => \n2_adj_1669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__36310\,
            in1 => \N__36136\,
            in2 => \N__36142\,
            in3 => \N__54613\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61833\,
            ce => \N__46427\,
            sr => \N__46350\
        );

    \mux_134_Mux_4_i4_3_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43084\,
            in1 => \N__54979\,
            in2 => \_gnd_net_\,
            in3 => \N__54415\,
            lcout => OPEN,
            ltout => \n4_adj_1670_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20463_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__54612\,
            in2 => \N__36139\,
            in3 => \N__51838\,
            lcout => n23402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20124_2_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38139\,
            in2 => \_gnd_net_\,
            in3 => \N__54413\,
            lcout => n22669,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_4_i1_3_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54414\,
            in1 => \_gnd_net_\,
            in2 => \N__44693\,
            in3 => \N__56096\,
            lcout => n1_adj_1668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10493_3_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36833\,
            in1 => \N__44677\,
            in2 => \_gnd_net_\,
            in3 => \N__46164\,
            lcout => n13219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__57176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36285\,
            lcout => \comm_spi.data_tx_7__N_871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62657\,
            in1 => \N__54024\,
            in2 => \_gnd_net_\,
            in3 => \N__38377\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__54809\,
            in1 => \N__62660\,
            in2 => \_gnd_net_\,
            in3 => \N__43555\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__54939\,
            in1 => \_gnd_net_\,
            in2 => \N__38488\,
            in3 => \N__62663\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i4_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__55071\,
            in1 => \N__62661\,
            in2 => \_gnd_net_\,
            in3 => \N__36262\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i5_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62658\,
            in1 => \N__55206\,
            in2 => \_gnd_net_\,
            in3 => \N__57919\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i6_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__53895\,
            in1 => \N__62662\,
            in2 => \_gnd_net_\,
            in3 => \N__36253\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \comm_buf_0__i7_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__62659\,
            in1 => \N__55937\,
            in2 => \N__36481\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61839\,
            ce => \N__61438\,
            sr => \N__64417\
        );

    \i16298_2_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36438\,
            lcout => n18996,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36400\,
            in1 => \N__62620\,
            in2 => \_gnd_net_\,
            in3 => \N__54025\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__62616\,
            in1 => \_gnd_net_\,
            in2 => \N__36394\,
            in3 => \N__54800\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41047\,
            in1 => \N__54940\,
            in2 => \_gnd_net_\,
            in3 => \N__62621\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62617\,
            in1 => \N__62789\,
            in2 => \_gnd_net_\,
            in3 => \N__36382\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55072\,
            in1 => \N__36373\,
            in2 => \_gnd_net_\,
            in3 => \N__62622\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62618\,
            in1 => \N__55207\,
            in2 => \_gnd_net_\,
            in3 => \N__36364\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53896\,
            in1 => \N__36355\,
            in2 => \_gnd_net_\,
            in3 => \N__62623\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_buf_2__i7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62619\,
            in1 => \_gnd_net_\,
            in2 => \N__55945\,
            in3 => \N__36727\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61844\,
            ce => \N__43462\,
            sr => \N__38425\
        );

    \comm_spi.data_tx_i2_12624_12625_set_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__37519\,
            in1 => \_gnd_net_\,
            in2 => \N__37573\,
            in3 => \N__37540\,
            lcout => \comm_spi.n15352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53697\,
            ce => 'H',
            sr => \N__36715\
        );

    \i4032_2_lut_3_lut_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__41019\,
            in1 => \N__38583\,
            in2 => \_gnd_net_\,
            in3 => \N__59367\,
            lcout => n6774,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i45_3_lut_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101110"
        )
    port map (
            in0 => \N__59364\,
            in1 => \N__61382\,
            in2 => \_gnd_net_\,
            in3 => \N__58652\,
            lcout => n40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_2_i111_3_lut_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38371\,
            in1 => \N__36630\,
            in2 => \_gnd_net_\,
            in3 => \N__59365\,
            lcout => OPEN,
            ltout => \n111_adj_1796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_2_i112_3_lut_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41066\,
            in2 => \N__36634\,
            in3 => \N__60597\,
            lcout => n112_adj_1797,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_2_i111_3_lut_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41067\,
            in1 => \N__36631\,
            in2 => \_gnd_net_\,
            in3 => \N__59366\,
            lcout => n111_adj_1750,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12640_12641_set_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36622\,
            in1 => \N__36598\,
            in2 => \_gnd_net_\,
            in3 => \N__36574\,
            lcout => \comm_spi.n15368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53698\,
            ce => 'H',
            sr => \N__36529\
        );

    \mux_125_Mux_5_i23_3_lut_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36501\,
            in1 => \N__59351\,
            in2 => \_gnd_net_\,
            in3 => \N__38821\,
            lcout => n23_adj_1773,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_7_i111_3_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59353\,
            in1 => \N__42376\,
            in2 => \_gnd_net_\,
            in3 => \N__38322\,
            lcout => n111_adj_1761,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_1_i111_3_lut_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41871\,
            in1 => \N__38391\,
            in2 => \_gnd_net_\,
            in3 => \N__59355\,
            lcout => n111_adj_1754,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_3_i16_3_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59352\,
            in1 => \N__36867\,
            in2 => \_gnd_net_\,
            in3 => \N__40069\,
            lcout => n16_adj_1738,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_4_i16_3_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49458\,
            in1 => \N__47268\,
            in2 => \_gnd_net_\,
            in3 => \N__59354\,
            lcout => n16_adj_1733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_51_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__37393\,
            in1 => \N__59446\,
            in2 => \N__56078\,
            in3 => \N__36841\,
            lcout => OPEN,
            ltout => \n11987_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__44714\,
            in1 => \N__38707\,
            in2 => \N__36817\,
            in3 => \N__43612\,
            lcout => \VAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61870\,
            ce => \N__36794\,
            sr => \N__37130\
        );

    \mux_125_Mux_4_i17_3_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37164\,
            in1 => \N__38792\,
            in2 => \_gnd_net_\,
            in3 => \N__59444\,
            lcout => n17_adj_1779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_258_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__59445\,
            in1 => \N__49146\,
            in2 => \N__43228\,
            in3 => \N__37392\,
            lcout => OPEN,
            ltout => \n11985_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__43933\,
            in1 => \N__37060\,
            in2 => \N__36802\,
            in3 => \N__43415\,
            lcout => \IAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61870\,
            ce => \N__36794\,
            sr => \N__37130\
        );

    \i1_2_lut_4_lut_adj_268_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__50890\,
            in1 => \N__55650\,
            in2 => \N__38758\,
            in3 => \N__37079\,
            lcout => n24_adj_1575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_269_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__50889\,
            in1 => \N__55649\,
            in2 => \N__38759\,
            in3 => \N__37037\,
            lcout => n24_adj_1601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_54_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__59363\,
            in1 => \N__45699\,
            in2 => \N__56582\,
            in3 => \N__37381\,
            lcout => n11984,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46842\,
            in1 => \N__50814\,
            in2 => \_gnd_net_\,
            in3 => \N__49848\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50815\,
            in1 => \N__48799\,
            in2 => \_gnd_net_\,
            in3 => \N__38215\,
            lcout => \buf_cfgRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_330_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40948\,
            in1 => \N__43872\,
            in2 => \_gnd_net_\,
            in3 => \N__39148\,
            lcout => acadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23438_bdd_4_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__37006\,
            in1 => \N__36997\,
            in2 => \N__36978\,
            in3 => \N__60072\,
            lcout => n23441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_5_i111_3_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36951\,
            in1 => \N__36933\,
            in2 => \_gnd_net_\,
            in3 => \N__59362\,
            lcout => OPEN,
            ltout => \n111_adj_1776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_5_i112_3_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36914\,
            in2 => \N__36883\,
            in3 => \N__60635\,
            lcout => n112_adj_1777,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_59_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__60636\,
            in1 => \_gnd_net_\,
            in2 => \N__60097\,
            in3 => \N__41020\,
            lcout => n11979,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i11_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39400\,
            in1 => \N__39799\,
            in2 => \N__44228\,
            in3 => \N__37284\,
            lcout => buf_adcdata_iac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37351\,
            in1 => \N__37333\,
            in2 => \N__41511\,
            in3 => \N__49844\,
            lcout => n24_adj_1513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_233_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__37315\,
            in1 => \N__37300\,
            in2 => \N__52743\,
            in3 => \N__37475\,
            lcout => n23_adj_1514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i20_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39798\,
            in1 => \N__37244\,
            in2 => \N__37285\,
            in3 => \N__37796\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57848\,
            in1 => \N__46852\,
            in2 => \N__40569\,
            in3 => \N__37476\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_0_i16_3_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37227\,
            in1 => \_gnd_net_\,
            in2 => \N__59513\,
            in3 => \N__47232\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i20_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39797\,
            in1 => \N__39401\,
            in2 => \N__37198\,
            in3 => \N__37163\,
            lcout => buf_adcdata_iac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47454\,
            in1 => \N__46846\,
            in2 => \_gnd_net_\,
            in3 => \N__39910\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__46845\,
            in1 => \N__57850\,
            in2 => \N__41510\,
            in3 => \N__46646\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i6_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57849\,
            in1 => \N__46738\,
            in2 => \N__40568\,
            in3 => \N__37486\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i2_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46736\,
            in1 => \N__47455\,
            in2 => \_gnd_net_\,
            in3 => \N__39927\,
            lcout => \SELIRNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_6_i23_3_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37485\,
            in1 => \N__59479\,
            in2 => \_gnd_net_\,
            in3 => \N__37477\,
            lcout => n23_adj_1767,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i4_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47356\,
            in1 => \N__46737\,
            in2 => \_gnd_net_\,
            in3 => \N__39875\,
            lcout => \VDC_RNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i1_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50540\,
            in1 => \N__50374\,
            in2 => \N__37447\,
            in3 => \N__42153\,
            lcout => \SIG_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61929\,
            ce => \N__42205\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i0_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50539\,
            in1 => \N__50373\,
            in2 => \N__40044\,
            in3 => \N__47233\,
            lcout => \SIG_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61929\,
            ce => \N__42205\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50372\,
            in1 => \N__50542\,
            in2 => \N__37414\,
            in3 => \N__40065\,
            lcout => \SIG_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61929\,
            ce => \N__42205\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i2_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50541\,
            in1 => \N__50375\,
            in2 => \N__37423\,
            in3 => \N__42358\,
            lcout => \SIG_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61929\,
            ce => \N__42205\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_12620_12621_reset_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37603\,
            in1 => \N__40288\,
            in2 => \_gnd_net_\,
            in3 => \N__37626\,
            lcout => \comm_spi.n15349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53568\,
            ce => 'H',
            sr => \N__37582\
        );

    \comm_spi.data_tx_i1_12620_12621_set_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__40287\,
            in2 => \_gnd_net_\,
            in3 => \N__37633\,
            lcout => \comm_spi.n15348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53588\,
            ce => 'H',
            sr => \N__37612\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37941\,
            lcout => \comm_spi.data_tx_7__N_860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43285\,
            in2 => \_gnd_net_\,
            in3 => \N__57116\,
            lcout => \comm_spi.data_tx_7__N_861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20218_4_lut_3_lut_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57117\,
            in1 => \N__37942\,
            in2 => \_gnd_net_\,
            in3 => \N__37556\,
            lcout => \comm_spi.n24037\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20449_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42520\,
            in1 => \N__54608\,
            in2 => \N__37921\,
            in3 => \N__51823\,
            lcout => n23390,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20253_4_lut_3_lut_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57114\,
            in1 => \N__43284\,
            in2 => \_gnd_net_\,
            in3 => \N__37598\,
            lcout => \comm_spi.n24040\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__37940\,
            in1 => \N__57113\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_12624_12625_reset_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37563\,
            in1 => \N__37533\,
            in2 => \_gnd_net_\,
            in3 => \N__37509\,
            lcout => \comm_spi.n15353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53601\,
            ce => 'H',
            sr => \N__40834\
        );

    \comm_spi.MISO_48_12606_12607_reset_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41970\,
            in1 => \N__42021\,
            in2 => \_gnd_net_\,
            in3 => \N__42003\,
            lcout => \comm_spi.n15335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12606_12607_resetC_net\,
            ce => 'H',
            sr => \N__40619\
        );

    \mux_134_Mux_1_i1_3_lut_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52121\,
            in1 => \N__44592\,
            in2 => \_gnd_net_\,
            in3 => \N__54372\,
            lcout => OPEN,
            ltout => \n1_adj_1674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__37909\,
            in1 => \N__37957\,
            in2 => \N__37945\,
            in3 => \N__54584\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61831\,
            ce => \N__46402\,
            sr => \N__46354\
        );

    \i19782_2_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40461\,
            in2 => \_gnd_net_\,
            in3 => \N__54370\,
            lcout => n22341,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_1_i2_3_lut_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41107\,
            in1 => \N__38307\,
            in2 => \_gnd_net_\,
            in3 => \N__54371\,
            lcout => n2_adj_1675,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_0_i19_3_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37903\,
            in1 => \N__37874\,
            in2 => \_gnd_net_\,
            in3 => \N__59436\,
            lcout => OPEN,
            ltout => \n19_adj_1590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_0_i22_3_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__38087\,
            in1 => \N__59993\,
            in2 => \N__37858\,
            in3 => \_gnd_net_\,
            lcout => n22_adj_1589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__59994\,
            in1 => \N__60467\,
            in2 => \N__46534\,
            in3 => \N__59437\,
            lcout => n21965,
            ltout => \n21965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_295_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57665\,
            in2 => \N__37843\,
            in3 => \N__63610\,
            lcout => n13093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i8_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37800\,
            in1 => \N__38117\,
            in2 => \N__38170\,
            in3 => \N__39810\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i4_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__38140\,
            in1 => \N__63611\,
            in2 => \N__55076\,
            in3 => \N__45562\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__39405\,
            in1 => \N__39758\,
            in2 => \N__38097\,
            in3 => \N__38118\,
            lcout => buf_adcdata_iac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_5_i19_3_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38071\,
            in1 => \N__38043\,
            in2 => \_gnd_net_\,
            in3 => \N__59435\,
            lcout => OPEN,
            ltout => \n19_adj_1729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20424_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__38017\,
            in1 => \N__59991\,
            in2 => \N__37993\,
            in3 => \N__60668\,
            lcout => n23354,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i6_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__37989\,
            in1 => \N__63612\,
            in2 => \N__53894\,
            in3 => \N__45569\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_3_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__59432\,
            in1 => \N__59992\,
            in2 => \_gnd_net_\,
            in3 => \N__60666\,
            lcout => n9_adj_1600,
            ltout => \n9_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4034_2_lut_3_lut_4_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__60667\,
            in1 => \N__41005\,
            in2 => \N__37975\,
            in3 => \N__59433\,
            lcout => n6776,
            ltout => \n6776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16190_3_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__45695\,
            in1 => \_gnd_net_\,
            in2 => \N__37972\,
            in3 => \N__45283\,
            lcout => n18890,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_1_i111_3_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43060\,
            in1 => \N__38395\,
            in2 => \_gnd_net_\,
            in3 => \N__59434\,
            lcout => n111_adj_1798,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_0_i127_3_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38521\,
            in1 => \N__61254\,
            in2 => \_gnd_net_\,
            in3 => \N__38530\,
            lcout => \comm_buf_0_7_N_543_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i16_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__57878\,
            in1 => \N__38472\,
            in2 => \N__43940\,
            in3 => \N__45401\,
            lcout => comm_test_buf_24_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i18_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45400\,
            in1 => \N__57879\,
            in2 => \N__40924\,
            in3 => \N__38367\,
            lcout => comm_test_buf_24_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16302_2_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60269\,
            in2 => \_gnd_net_\,
            in3 => \N__58855\,
            lcout => n112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_7_i111_3_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58857\,
            in1 => \N__38353\,
            in2 => \_gnd_net_\,
            in3 => \N__38329\,
            lcout => n111_adj_1719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10475_3_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38297\,
            in1 => \N__44565\,
            in2 => \_gnd_net_\,
            in3 => \N__46195\,
            lcout => n13201,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20538_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__58856\,
            in1 => \N__38266\,
            in2 => \N__60397\,
            in3 => \N__38233\,
            lcout => n23486,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19795_2_lut_3_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__38582\,
            in1 => \N__60980\,
            in2 => \_gnd_net_\,
            in3 => \N__58648\,
            lcout => n22354,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_12612_12613_set_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38191\,
            in1 => \N__41980\,
            in2 => \_gnd_net_\,
            in3 => \N__38443\,
            lcout => \comm_spi.n15340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12612_12613_setC_net\,
            ce => 'H',
            sr => \N__41914\
        );

    \i16457_2_lut_3_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__62610\,
            in1 => \N__40890\,
            in2 => \_gnd_net_\,
            in3 => \N__63990\,
            lcout => n14_adj_1655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16462_2_lut_3_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__63991\,
            in1 => \N__43914\,
            in2 => \_gnd_net_\,
            in3 => \N__62611\,
            lcout => n14_adj_1608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__62609\,
            in1 => \N__63988\,
            in2 => \_gnd_net_\,
            in3 => \N__51614\,
            lcout => n11254,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_193_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__63989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63603\,
            lcout => n21968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12520_2_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__63604\,
            in1 => \_gnd_net_\,
            in2 => \N__62676\,
            in3 => \_gnd_net_\,
            lcout => n15238,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12773_2_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63606\,
            in2 => \_gnd_net_\,
            in3 => \N__43458\,
            lcout => n15496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12780_2_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__63605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41031\,
            lcout => n15503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19343_4_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__60595\,
            in1 => \N__59321\,
            in2 => \N__38416\,
            in3 => \N__46864\,
            lcout => OPEN,
            ltout => \n22270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_20503_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__59995\,
            in1 => \N__38500\,
            in2 => \N__38398\,
            in3 => \N__60992\,
            lcout => OPEN,
            ltout => \n23450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23450_bdd_4_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__60993\,
            in1 => \N__43474\,
            in2 => \N__38545\,
            in3 => \N__38542\,
            lcout => n23453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_0_i112_3_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48993\,
            in1 => \N__38458\,
            in2 => \_gnd_net_\,
            in3 => \N__60596\,
            lcout => n112_adj_1583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23522_bdd_4_lut_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__38512\,
            in1 => \N__60594\,
            in2 => \N__52642\,
            in3 => \N__44116\,
            lcout => n22267,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_2_i127_3_lut_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38494\,
            in1 => \N__61253\,
            in2 => \_gnd_net_\,
            in3 => \N__41413\,
            lcout => \comm_buf_0_7_N_543_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_0_i111_3_lut_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59320\,
            in1 => \N__38476\,
            in2 => \_gnd_net_\,
            in3 => \N__48957\,
            lcout => n111_adj_1584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_254_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44336\,
            in1 => \N__51985\,
            in2 => \N__51948\,
            in3 => \N__49819\,
            lcout => n20_adj_1804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51352\,
            in1 => \N__51944\,
            in2 => \_gnd_net_\,
            in3 => \N__47112\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39192\,
            in1 => \N__47424\,
            in2 => \_gnd_net_\,
            in3 => \N__51353\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_253_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__50128\,
            in1 => \N__50086\,
            in2 => \N__38690\,
            in3 => \N__39191\,
            lcout => n21_adj_1803,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38694\,
            in1 => \N__47363\,
            in2 => \_gnd_net_\,
            in3 => \N__51354\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20478_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__38661\,
            in1 => \N__60631\,
            in2 => \N__38619\,
            in3 => \N__59305\,
            lcout => n23348,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19165_3_lut_1_lut_2_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41015\,
            in2 => \_gnd_net_\,
            in3 => \N__38584\,
            lcout => n22092,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_331_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44613\,
            in1 => \N__43865\,
            in2 => \_gnd_net_\,
            in3 => \N__38866\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_2_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47815\,
            in1 => \N__47814\,
            in2 => \N__47769\,
            in3 => \N__38560\,
            lcout => n7,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => n20652,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_3_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__40204\,
            in1 => \N__40203\,
            in2 => \N__47773\,
            in3 => \N__38557\,
            lcout => n7_adj_1629,
            ltout => OPEN,
            carryin => n20652,
            carryout => n20653,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_4_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41790\,
            in1 => \N__41789\,
            in2 => \N__47770\,
            in3 => \N__38554\,
            lcout => n7_adj_1627,
            ltout => OPEN,
            carryin => n20653,
            carryout => n20654,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_5_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41625\,
            in1 => \N__41624\,
            in2 => \N__47774\,
            in3 => \N__38551\,
            lcout => n7_adj_1626,
            ltout => OPEN,
            carryin => n20654,
            carryout => n20655,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_6_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__44164\,
            in1 => \N__44163\,
            in2 => \N__47771\,
            in3 => \N__38548\,
            lcout => n7_adj_1624,
            ltout => OPEN,
            carryin => n20655,
            carryout => n20656,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_7_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__56503\,
            in1 => \N__56502\,
            in2 => \N__47776\,
            in3 => \N__38887\,
            lcout => n7_adj_1622,
            ltout => OPEN,
            carryin => n20656,
            carryout => n20657,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_8_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45148\,
            in1 => \N__45147\,
            in2 => \N__47772\,
            in3 => \N__38884\,
            lcout => n7_adj_1620,
            ltout => OPEN,
            carryin => n20657,
            carryout => n20658,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_9_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45007\,
            in1 => \N__45006\,
            in2 => \N__47775\,
            in3 => \N__38881\,
            lcout => n7_adj_1618,
            ltout => OPEN,
            carryin => n20658,
            carryout => n20659,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_10_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__44953\,
            in1 => \N__44952\,
            in2 => \N__47784\,
            in3 => \N__38878\,
            lcout => n7_adj_1616,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => n20660,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_122_11_lut_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42332\,
            in1 => \N__42333\,
            in2 => \N__47783\,
            in3 => \N__38875\,
            lcout => n7_adj_1614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20523_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__59438\,
            in1 => \N__38871\,
            in2 => \N__60663\,
            in3 => \N__44080\,
            lcout => n23480,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_58_i14_2_lut_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38839\,
            in2 => \_gnd_net_\,
            in3 => \N__38816\,
            lcout => n14_adj_1599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__38817\,
            in1 => \_gnd_net_\,
            in2 => \N__55283\,
            in3 => \N__46819\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_121_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__38793\,
            in1 => \N__55640\,
            in2 => \N__38773\,
            in3 => \N__50891\,
            lcout => n24_adj_1505,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16164_3_lut_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49293\,
            in1 => \N__41626\,
            in2 => \_gnd_net_\,
            in3 => \N__56469\,
            lcout => n18865,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19240_3_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39196\,
            in1 => \N__39133\,
            in2 => \_gnd_net_\,
            in3 => \N__59439\,
            lcout => n22167,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_3_i15_4_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__41652\,
            in1 => \N__63607\,
            in2 => \N__57746\,
            in3 => \N__41641\,
            lcout => \data_index_9_N_236_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_232_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38983\,
            in1 => \N__38965\,
            in2 => \N__52811\,
            in3 => \N__55469\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__55470\,
            in1 => \N__47517\,
            in2 => \N__46844\,
            in3 => \_gnd_net_\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__56839\,
            in1 => \_gnd_net_\,
            in2 => \N__46843\,
            in3 => \N__52742\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_234_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__38947\,
            in1 => \N__38929\,
            in2 => \N__39855\,
            in3 => \N__39908\,
            lcout => OPEN,
            ltout => \n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_238_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38911\,
            in1 => \N__38902\,
            in2 => \N__38896\,
            in3 => \N__38893\,
            lcout => n30_adj_1743,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47367\,
            in2 => \N__39856\,
            in3 => \N__46810\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61916\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16464_2_lut_3_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__63992\,
            in1 => \N__49232\,
            in2 => \_gnd_net_\,
            in3 => \N__62692\,
            lcout => n14_adj_1610,
            ltout => \n14_adj_1610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__49683\,
            in1 => \_gnd_net_\,
            in2 => \N__39985\,
            in3 => \N__46847\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_240_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__39981\,
            in1 => \N__49682\,
            in2 => \N__39964\,
            in3 => \N__47030\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19239_3_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39926\,
            in1 => \N__59441\,
            in2 => \_gnd_net_\,
            in3 => \N__39909\,
            lcout => n22166,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_4_i23_3_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__59440\,
            in1 => \_gnd_net_\,
            in2 => \N__39879\,
            in3 => \N__39854\,
            lcout => n23_adj_1783,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__47031\,
            in1 => \N__57856\,
            in2 => \N__49142\,
            in3 => \N__46848\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i9_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__39806\,
            in1 => \N__39385\,
            in2 => \N__39223\,
            in3 => \N__52704\,
            lcout => buf_adcdata_iac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i1_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__50737\,
            in1 => \N__52091\,
            in2 => \N__57880\,
            in3 => \N__42152\,
            lcout => buf_dds0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__40171\,
            in1 => \N__40180\,
            in2 => \N__57871\,
            in3 => \N__63609\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i8_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50736\,
            in1 => \N__48857\,
            in2 => \_gnd_net_\,
            in3 => \N__40226\,
            lcout => buf_dds0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6651_3_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52090\,
            in1 => \N__40196\,
            in2 => \_gnd_net_\,
            in3 => \N__56474\,
            lcout => n8_adj_1630,
            ltout => \n8_adj_1630_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_1_i15_4_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__63608\,
            in1 => \N__57833\,
            in2 => \N__40174\,
            in3 => \N__40170\,
            lcout => \data_index_9_N_236_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i3_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57834\,
            in1 => \N__50738\,
            in2 => \N__49311\,
            in3 => \N__40064\,
            lcout => buf_dds0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i3_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__56849\,
            in1 => \N__46750\,
            in2 => \_gnd_net_\,
            in3 => \N__52763\,
            lcout => \SELIRNG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.MOSI_31_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40045\,
            in1 => \N__40011\,
            in2 => \_gnd_net_\,
            in3 => \N__50368\,
            lcout => \DDS_MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61970\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12598_12599_set_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42498\,
            lcout => \comm_spi.n15326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61824\,
            ce => 'H',
            sr => \N__42166\
        );

    \comm_spi.i20203_4_lut_3_lut_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42499\,
            in1 => \N__40000\,
            in2 => \_gnd_net_\,
            in3 => \N__57130\,
            lcout => \comm_spi.n24016\,
            ltout => \comm_spi.n24016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12600_3_lut_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39994\,
            in1 => \_gnd_net_\,
            in2 => \N__39988\,
            in3 => \N__42766\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12594_12595_set_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__64676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n15322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53617\,
            ce => 'H',
            sr => \N__40276\
        );

    \secclk_cnt_3785_3786__i1_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45223\,
            in2 => \_gnd_net_\,
            in3 => \N__40264\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => n20790,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42405\,
            in2 => \_gnd_net_\,
            in3 => \N__40261\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n20790,
            carryout => n20791,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42865\,
            in2 => \_gnd_net_\,
            in3 => \N__40258\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n20791,
            carryout => n20792,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42922\,
            in2 => \_gnd_net_\,
            in3 => \N__40255\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n20792,
            carryout => n20793,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45168\,
            in2 => \_gnd_net_\,
            in3 => \N__40252\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n20793,
            carryout => n20794,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42391\,
            in2 => \_gnd_net_\,
            in3 => \N__40249\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n20794,
            carryout => n20795,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42961\,
            in2 => \_gnd_net_\,
            in3 => \N__40246\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n20795,
            carryout => n20796,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42892\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n20796,
            carryout => n20797,
            clk => \N__48400\,
            ce => 'H',
            sr => \N__42846\
        );

    \secclk_cnt_3785_3786__i9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42418\,
            in2 => \_gnd_net_\,
            in3 => \N__40315\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => n20798,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42994\,
            in2 => \_gnd_net_\,
            in3 => \N__40312\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n20798,
            carryout => n20799,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42936\,
            in2 => \_gnd_net_\,
            in3 => \N__40309\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n20799,
            carryout => n20800,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i12_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45183\,
            in2 => \_gnd_net_\,
            in3 => \N__40306\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n20800,
            carryout => n20801,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i13_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40341\,
            in2 => \_gnd_net_\,
            in3 => \N__40303\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n20801,
            carryout => n20802,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i14_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42879\,
            in2 => \_gnd_net_\,
            in3 => \N__40300\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n20802,
            carryout => n20803,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i15_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42949\,
            in2 => \_gnd_net_\,
            in3 => \N__40297\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n20803,
            carryout => n20804,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i16_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42430\,
            in2 => \_gnd_net_\,
            in3 => \N__40294\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n20804,
            carryout => n20805,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__42845\
        );

    \secclk_cnt_3785_3786__i17_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42904\,
            in2 => \_gnd_net_\,
            in3 => \N__40291\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => n20806,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i18_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42981\,
            in2 => \_gnd_net_\,
            in3 => \N__40387\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n20806,
            carryout => n20807,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i19_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45207\,
            in2 => \_gnd_net_\,
            in3 => \N__40384\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n20807,
            carryout => n20808,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i20_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40369\,
            in2 => \_gnd_net_\,
            in3 => \N__40381\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n20808,
            carryout => n20809,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i21_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43018\,
            in2 => \_gnd_net_\,
            in3 => \N__40378\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n20809,
            carryout => n20810,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i22_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40357\,
            in2 => \_gnd_net_\,
            in3 => \N__40375\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n20810,
            carryout => n20811,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \secclk_cnt_3785_3786__i23_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40327\,
            in2 => \_gnd_net_\,
            in3 => \N__40372\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48403\,
            ce => 'H',
            sr => \N__42847\
        );

    \i6_4_lut_adj_204_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40368\,
            in1 => \N__40356\,
            in2 => \N__40345\,
            in3 => \N__40326\,
            lcout => n14_adj_1678,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_287_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__63483\,
            in1 => \N__63163\,
            in2 => \N__64101\,
            in3 => \N__51542\,
            lcout => n15378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_333_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__63162\,
            in1 => \N__64090\,
            in2 => \N__51546\,
            in3 => \N__63482\,
            lcout => n13076,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16454_2_lut_3_lut_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__64091\,
            in1 => \N__40563\,
            in2 => \_gnd_net_\,
            in3 => \N__62624\,
            lcout => n14_adj_1652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__40465\,
            in1 => \N__63484\,
            in2 => \N__54823\,
            in3 => \N__45570\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_127_Mux_2_i30_3_lut_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40450\,
            in1 => \N__40438\,
            in2 => \_gnd_net_\,
            in3 => \N__60991\,
            lcout => n30_adj_1708,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_215_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__63485\,
            in1 => \N__64095\,
            in2 => \N__63189\,
            in3 => \N__56884\,
            lcout => n12585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i13_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__57764\,
            in1 => \N__55529\,
            in2 => \N__45339\,
            in3 => \N__50688\,
            lcout => buf_dds0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i2_3_lut_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40424\,
            in1 => \N__40783\,
            in2 => \_gnd_net_\,
            in3 => \N__54407\,
            lcout => n2_adj_1663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19758_2_lut_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__54408\,
            in1 => \N__43071\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n22331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20429_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__40669\,
            in1 => \N__54599\,
            in2 => \N__40399\,
            in3 => \N__51822\,
            lcout => OPEN,
            ltout => \n23360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__54600\,
            in1 => \N__40663\,
            in2 => \N__40396\,
            in3 => \N__40393\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61842\,
            ce => \N__46403\,
            sr => \N__46351\
        );

    \mux_134_Mux_7_i4_3_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__53908\,
            in1 => \N__43147\,
            in2 => \_gnd_net_\,
            in3 => \N__54405\,
            lcout => n4_adj_1664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i1_3_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54406\,
            in1 => \N__46622\,
            in2 => \_gnd_net_\,
            in3 => \N__55841\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20213_4_lut_3_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41963\,
            in1 => \N__40643\,
            in2 => \_gnd_net_\,
            in3 => \N__57111\,
            lcout => \comm_spi.n15333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__57112\,
            in1 => \_gnd_net_\,
            in2 => \N__40650\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_862\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_2_i4_3_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43354\,
            in1 => \N__54838\,
            in2 => \_gnd_net_\,
            in3 => \N__54398\,
            lcout => n4_adj_1673,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19747_2_lut_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__54399\,
            in1 => \_gnd_net_\,
            in2 => \N__45517\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n22342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20454_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__40597\,
            in1 => \N__54601\,
            in2 => \N__40591\,
            in3 => \N__51830\,
            lcout => n23396,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_2_i1_3_lut_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54401\,
            in1 => \_gnd_net_\,
            in2 => \N__40939\,
            in3 => \N__52926\,
            lcout => OPEN,
            ltout => \n1_adj_1671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__40588\,
            in1 => \N__54602\,
            in2 => \N__40582\,
            in3 => \N__40579\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61848\,
            ce => \N__46431\,
            sr => \N__46349\
        );

    \mux_134_Mux_2_i2_3_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54400\,
            in1 => \N__41128\,
            in2 => \_gnd_net_\,
            in3 => \N__40973\,
            lcout => n2_adj_1672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10481_3_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40974\,
            in1 => \N__40925\,
            in2 => \_gnd_net_\,
            in3 => \N__46163\,
            lcout => n13207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__57110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40845\,
            lcout => \comm_spi.data_tx_7__N_877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__54016\,
            in1 => \N__40816\,
            in2 => \_gnd_net_\,
            in3 => \N__62653\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62652\,
            in1 => \_gnd_net_\,
            in2 => \N__55936\,
            in3 => \N__40801\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i6_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53879\,
            in1 => \N__40774\,
            in2 => \_gnd_net_\,
            in3 => \N__62656\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i5_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62648\,
            in1 => \_gnd_net_\,
            in2 => \N__55194\,
            in3 => \N__40738\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i4_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55077\,
            in1 => \N__40717\,
            in2 => \_gnd_net_\,
            in3 => \N__62655\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i3_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62647\,
            in1 => \N__62790\,
            in2 => \_gnd_net_\,
            in3 => \N__40687\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i2_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__54938\,
            in1 => \N__41143\,
            in2 => \_gnd_net_\,
            in3 => \N__62654\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \comm_buf_3__i1_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__54816\,
            in1 => \_gnd_net_\,
            in2 => \N__62685\,
            in3 => \N__41122\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61855\,
            ce => \N__41038\,
            sr => \N__41095\
        );

    \mux_127_Mux_2_i127_3_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41080\,
            in1 => \N__41071\,
            in2 => \_gnd_net_\,
            in3 => \N__61182\,
            lcout => \comm_buf_2_7_N_575_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_316_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__54136\,
            in1 => \N__54085\,
            in2 => \_gnd_net_\,
            in3 => \N__48889\,
            lcout => n12880,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__45933\,
            in1 => \N__45995\,
            in2 => \N__53893\,
            in3 => \N__61183\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__58585\,
            in1 => \N__58469\,
            in2 => \N__61260\,
            in3 => \N__60793\,
            lcout => n21886,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_310_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__60792\,
            in1 => \N__61178\,
            in2 => \N__58491\,
            in3 => \N__58584\,
            lcout => n12,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58836\,
            in2 => \N__40981\,
            in3 => \_gnd_net_\,
            lcout => n12015,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_338_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__59672\,
            in1 => \N__41349\,
            in2 => \N__63075\,
            in3 => \N__41400\,
            lcout => n11258,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12830_2_lut_3_lut_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64089\,
            in2 => \N__44040\,
            in3 => \N__62615\,
            lcout => n15553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16466_2_lut_3_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__52909\,
            in1 => \N__62689\,
            in2 => \_gnd_net_\,
            in3 => \N__64088\,
            lcout => n14_adj_1612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23288_bdd_4_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__43660\,
            in1 => \N__41326\,
            in2 => \N__41311\,
            in3 => \N__59999\,
            lcout => n23291,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__60000\,
            in1 => \N__63078\,
            in2 => \N__41266\,
            in3 => \N__60468\,
            lcout => n9324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51348\,
            in1 => \_gnd_net_\,
            in2 => \N__48941\,
            in3 => \N__44340\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_372_i8_2_lut_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__60469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60001\,
            lcout => OPEN,
            ltout => \n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_210_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__41265\,
            in1 => \N__63726\,
            in2 => \N__41254\,
            in3 => \N__63079\,
            lcout => n11172,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_3_i19_3_lut_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41251\,
            in1 => \N__41220\,
            in2 => \_gnd_net_\,
            in3 => \N__59306\,
            lcout => n19_adj_1739,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_73_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__63081\,
            in1 => \N__41194\,
            in2 => \N__57844\,
            in3 => \N__63725\,
            lcout => n13211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__41164\,
            in1 => \N__41533\,
            in2 => \N__44296\,
            in3 => \N__51917\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_7_i23_3_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46024\,
            in1 => \N__59307\,
            in2 => \_gnd_net_\,
            in3 => \N__41512\,
            lcout => n23_adj_1756,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_313_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51685\,
            in1 => \N__41470\,
            in2 => \N__44092\,
            in3 => \N__43573\,
            lcout => n30_adj_1769,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23546_bdd_4_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__41455\,
            in1 => \N__60002\,
            in2 => \N__41446\,
            in3 => \N__44140\,
            lcout => OPEN,
            ltout => \n23549_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19247_3_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41431\,
            in2 => \N__41416\,
            in3 => \N__60994\,
            lcout => n22174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44134\,
            in1 => \N__61348\,
            in2 => \_gnd_net_\,
            in3 => \N__41407\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61903\,
            ce => \N__46678\,
            sr => \N__48291\
        );

    \comm_length_i1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__61347\,
            in1 => \N__41389\,
            in2 => \_gnd_net_\,
            in3 => \N__60664\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61903\,
            ce => \N__46678\,
            sr => \N__48291\
        );

    \i1_2_lut_adj_244_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43818\,
            in2 => \_gnd_net_\,
            in3 => \N__41544\,
            lcout => n17650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_331_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63080\,
            in2 => \_gnd_net_\,
            in3 => \N__41353\,
            lcout => n21983,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20055_2_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41806\,
            in2 => \_gnd_net_\,
            in3 => \N__59322\,
            lcout => n22301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63735\,
            in1 => \N__41773\,
            in2 => \N__57778\,
            in3 => \N__41764\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6641_3_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52888\,
            in1 => \N__41791\,
            in2 => \_gnd_net_\,
            in3 => \N__56462\,
            lcout => n8_adj_1628,
            ltout => \n8_adj_1628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_2_i15_4_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57692\,
            in1 => \N__63618\,
            in2 => \N__41767\,
            in3 => \N__41763\,
            lcout => \data_index_9_N_236_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__52889\,
            in1 => \N__46818\,
            in2 => \N__52816\,
            in3 => \N__57700\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63736\,
            in1 => \N__41653\,
            in2 => \N__57779\,
            in3 => \N__41640\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_236_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__41608\,
            in1 => \N__44105\,
            in2 => \N__41587\,
            in3 => \N__41575\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_241_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43972\,
            in1 => \N__41569\,
            in2 => \N__41560\,
            in3 => \N__41557\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_321_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__51380\,
            in1 => \N__46486\,
            in2 => \N__63723\,
            in3 => \N__57693\,
            lcout => n13141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_1_i16_3_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42154\,
            in1 => \N__42132\,
            in2 => \_gnd_net_\,
            in3 => \N__59442\,
            lcout => n16_adj_1751,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_2_i16_3_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42103\,
            in1 => \N__42350\,
            in2 => \_gnd_net_\,
            in3 => \N__59443\,
            lcout => OPEN,
            ltout => \n16_adj_1746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19221_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42069\,
            in2 => \N__42034\,
            in3 => \N__60599\,
            lcout => n22148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_12606_12607_set_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42031\,
            in1 => \N__42007\,
            in2 => \_gnd_net_\,
            in3 => \N__41985\,
            lcout => \comm_spi.n15334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12606_12607_setC_net\,
            ce => 'H',
            sr => \N__41913\
        );

    \mux_125_Mux_1_i112_3_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41872\,
            in1 => \N__41836\,
            in2 => \_gnd_net_\,
            in3 => \N__60598\,
            lcout => n112_adj_1799,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4594_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49129\,
            in1 => \N__47813\,
            in2 => \_gnd_net_\,
            in3 => \N__56458\,
            lcout => n8_adj_1605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_207_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__41824\,
            in1 => \N__63194\,
            in2 => \N__63784\,
            in3 => \N__57703\,
            lcout => OPEN,
            ltout => \n12056_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds0_307_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__57705\,
            in1 => \N__47575\,
            in2 => \N__41809\,
            in3 => \N__63777\,
            lcout => trig_dds0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i4_4_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__47662\,
            in1 => \N__44737\,
            in2 => \N__44763\,
            in3 => \N__50614\,
            lcout => \SIG_DDS.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i23_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__42372\,
            in1 => \N__46647\,
            in2 => \N__45427\,
            in3 => \N__57706\,
            lcout => comm_test_buf_24_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i2_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57704\,
            in1 => \N__50776\,
            in2 => \N__52925\,
            in3 => \N__42351\,
            lcout => buf_dds0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6591_3_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__56459\,
            in1 => \_gnd_net_\,
            in2 => \N__55837\,
            in3 => \N__44999\,
            lcout => n8_adj_1619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6571_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44632\,
            in1 => \N__42334\,
            in2 => \_gnd_net_\,
            in3 => \N__56460\,
            lcout => n8_adj_1615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6581_3_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__56461\,
            in1 => \N__43947\,
            in2 => \_gnd_net_\,
            in3 => \N__44940\,
            lcout => n8_adj_1617,
            ltout => \n8_adj_1617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_8_i15_4_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57702\,
            in1 => \N__63724\,
            in2 => \N__42301\,
            in3 => \N__44970\,
            lcout => \data_index_9_N_236_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i2_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50460\,
            in2 => \_gnd_net_\,
            in3 => \N__50364\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61983\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i20129_4_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000110"
        )
    port map (
            in0 => \N__50592\,
            in1 => \N__50459\,
            in2 => \N__47584\,
            in3 => \N__50363\,
            lcout => \SIG_DDS.n13338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57118\,
            lcout => \comm_spi.iclk_N_850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12602_12603_reset_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n15331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61825\,
            ce => 'H',
            sr => \N__44794\
        );

    \comm_spi.iclk_40_12598_12599_reset_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42490\,
            lcout => \comm_spi.n15327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61827\,
            ce => 'H',
            sr => \N__42442\
        );

    \comm_spi.data_rx_i0_12616_12617_reset_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47959\,
            in1 => \N__44785\,
            in2 => \_gnd_net_\,
            in3 => \N__45459\,
            lcout => \comm_spi.n15345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53634\,
            ce => 'H',
            sr => \N__42511\
        );

    \ADC_VDC.genclk.t_clk_24_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64227\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VDC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t_clk_24C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_1_i4_3_lut_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43333\,
            in1 => \N__54709\,
            in2 => \_gnd_net_\,
            in3 => \N__54409\,
            lcout => n4_adj_1676,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__57121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47542\,
            lcout => \comm_spi.DOUT_7__N_835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__42491\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57120\,
            lcout => \comm_spi.iclk_N_851\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42429\,
            in1 => \N__42417\,
            in2 => \N__42406\,
            in3 => \N__42390\,
            lcout => OPEN,
            ltout => \n25_adj_1717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_205_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45154\,
            in1 => \N__42853\,
            in2 => \N__42379\,
            in3 => \N__42910\,
            lcout => OPEN,
            ltout => \n20922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__42967\,
            in1 => \N__43017\,
            in2 => \N__43006\,
            in3 => \N__43003\,
            lcout => n15420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42993\,
            in2 => \_gnd_net_\,
            in3 => \N__42982\,
            lcout => n10_adj_1679,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_203_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42960\,
            in1 => \N__42948\,
            in2 => \N__42937\,
            in3 => \N__42921\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42903\,
            in1 => \N__42891\,
            in2 => \N__42880\,
            in3 => \N__42864\,
            lcout => n26_adj_1715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SecClk_295_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42792\,
            in2 => \_gnd_net_\,
            in3 => \N__42826\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_374_i9_2_lut_3_lut_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__59189\,
            in1 => \N__59969\,
            in2 => \_gnd_net_\,
            in3 => \N__60498\,
            lcout => n9_adj_1596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9640_1_lut_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52658\,
            lcout => n12366,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19311_3_lut_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__58204\,
            in1 => \N__62637\,
            in2 => \_gnd_net_\,
            in3 => \N__63082\,
            lcout => n22238,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i7_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__43072\,
            in1 => \N__63487\,
            in2 => \N__55941\,
            in3 => \N__45558\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_test_buf_24_i17_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__57520\,
            in1 => \N__43056\,
            in2 => \N__44631\,
            in3 => \N__45372\,
            lcout => comm_test_buf_24_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__51165\,
            in1 => \N__55935\,
            in2 => \N__45955\,
            in3 => \N__45977\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__63489\,
            in1 => \N__53990\,
            in2 => \N__43042\,
            in3 => \N__45557\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12808_3_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__46390\,
            in1 => \N__63486\,
            in2 => \_gnd_net_\,
            in3 => \N__51164\,
            lcout => n15531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i5_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__45556\,
            in1 => \N__45714\,
            in2 => \N__55193\,
            in3 => \N__63490\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16114_3_lut_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43041\,
            in1 => \N__43226\,
            in2 => \_gnd_net_\,
            in3 => \N__54588\,
            lcout => n18816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16116_3_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54587\,
            in1 => \N__43171\,
            in2 => \_gnd_net_\,
            in3 => \N__49122\,
            lcout => OPEN,
            ltout => \n18818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20434_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__43240\,
            in1 => \N__54362\,
            in2 => \N__43024\,
            in3 => \N__51821\,
            lcout => OPEN,
            ltout => \n23372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i0_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__54363\,
            in1 => \N__43234\,
            in2 => \N__43021\,
            in3 => \N__43294\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61849\,
            ce => \N__46404\,
            sr => \N__46352\
        );

    \i19938_2_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43249\,
            in2 => \_gnd_net_\,
            in3 => \N__54586\,
            lcout => n22338,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16113_3_lut_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54589\,
            in1 => \_gnd_net_\,
            in2 => \N__43956\,
            in3 => \N__53938\,
            lcout => n18815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16121_3_lut_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43227\,
            in1 => \N__43948\,
            in2 => \_gnd_net_\,
            in3 => \N__46201\,
            lcout => n18823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43186\,
            in1 => \N__62629\,
            in2 => \_gnd_net_\,
            in3 => \N__54015\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i7_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62628\,
            in1 => \_gnd_net_\,
            in2 => \N__55931\,
            in3 => \N__43165\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i6_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53856\,
            in1 => \N__43141\,
            in2 => \_gnd_net_\,
            in3 => \N__62632\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i5_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62627\,
            in1 => \N__55160\,
            in2 => \_gnd_net_\,
            in3 => \N__43114\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i4_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55067\,
            in1 => \N__43099\,
            in2 => \_gnd_net_\,
            in3 => \N__62631\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i3_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62626\,
            in1 => \_gnd_net_\,
            in2 => \N__62779\,
            in3 => \N__43387\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i2_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__54931\,
            in1 => \N__43369\,
            in2 => \_gnd_net_\,
            in3 => \N__62630\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_buf_5__i1_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62625\,
            in1 => \N__54788\,
            in2 => \_gnd_net_\,
            in3 => \N__43348\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61856\,
            ce => \N__45886\,
            sr => \N__45736\
        );

    \comm_cmd_i0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__58844\,
            in1 => \N__54020\,
            in2 => \N__45953\,
            in3 => \N__45996\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__59703\,
            in1 => \N__45998\,
            in2 => \N__45954\,
            in3 => \N__54930\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__45942\,
            in1 => \N__45997\,
            in2 => \N__62794\,
            in3 => \N__60865\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_188_i9_2_lut_3_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__59702\,
            in1 => \N__60248\,
            in2 => \_gnd_net_\,
            in3 => \N__58842\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_60_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__61231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58614\,
            lcout => n8_adj_1504,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_20553_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__48706\,
            in1 => \N__60249\,
            in2 => \N__43321\,
            in3 => \N__58843\,
            lcout => OPEN,
            ltout => \n23504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23504_bdd_4_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__60250\,
            in1 => \N__43543\,
            in2 => \N__43519\,
            in3 => \N__43509\,
            lcout => n22288,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i1_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57620\,
            in1 => \N__46749\,
            in2 => \N__44617\,
            in3 => \N__49866\,
            lcout => \DDS_RNG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_315_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__63045\,
            in1 => \N__61300\,
            in2 => \N__43650\,
            in3 => \N__58608\,
            lcout => n21964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_309_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__54081\,
            in1 => \N__63046\,
            in2 => \N__54161\,
            in3 => \N__45865\,
            lcout => n12838,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20382_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__45829\,
            in1 => \N__60262\,
            in2 => \N__49012\,
            in3 => \N__59812\,
            lcout => n23306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19135_2_lut_3_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__58609\,
            in1 => \N__58365\,
            in2 => \_gnd_net_\,
            in3 => \N__61232\,
            lcout => n22061,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__58483\,
            in1 => \N__45941\,
            in2 => \N__55081\,
            in3 => \N__46008\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_374_i10_2_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58482\,
            in2 => \_gnd_net_\,
            in3 => \N__60879\,
            lcout => n6,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_62_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__43435\,
            in1 => \N__43633\,
            in2 => \N__43426\,
            in3 => \N__46481\,
            lcout => n21938,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__45940\,
            in1 => \N__58615\,
            in2 => \N__46012\,
            in3 => \N__55189\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20372_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__59822\,
            in1 => \N__43699\,
            in2 => \N__43687\,
            in3 => \N__60353\,
            lcout => n23288,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__46849\,
            in1 => \N__57619\,
            in2 => \N__51925\,
            in3 => \N__56577\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57618\,
            in1 => \N__46850\,
            in2 => \N__52142\,
            in3 => \N__52233\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51362\,
            in1 => \_gnd_net_\,
            in2 => \N__52842\,
            in3 => \N__47154\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61888\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19814_3_lut_4_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__61267\,
            in1 => \N__60880\,
            in2 => \N__59973\,
            in3 => \N__58607\,
            lcout => OPEN,
            ltout => \n22396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19906_4_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__60352\,
            in1 => \N__56170\,
            in2 => \N__43654\,
            in3 => \N__58487\,
            lcout => n22397,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_56_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001111"
        )
    port map (
            in0 => \N__61268\,
            in1 => \N__46453\,
            in2 => \N__43651\,
            in3 => \N__43632\,
            lcout => n21929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_250_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__55490\,
            in1 => \N__54658\,
            in2 => \N__52405\,
            in3 => \N__52832\,
            lcout => n22_adj_1801,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_1_i127_3_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43567\,
            in1 => \N__61291\,
            in2 => \_gnd_net_\,
            in3 => \N__50965\,
            lcout => \comm_buf_0_7_N_543_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_255_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__52482\,
            in1 => \N__52549\,
            in2 => \N__52206\,
            in3 => \N__52258\,
            lcout => n18_adj_1699,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__52205\,
            in1 => \N__47185\,
            in2 => \N__51338\,
            in3 => \_gnd_net_\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_302_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__46203\,
            in1 => \N__63051\,
            in2 => \N__63762\,
            in3 => \N__57610\,
            lcout => n13257,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47515\,
            in2 => \N__55497\,
            in3 => \N__51310\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_235_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44017\,
            in1 => \N__52505\,
            in2 => \N__43996\,
            in3 => \N__52229\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_332_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43960\,
            in1 => \N__43873\,
            in2 => \_gnd_net_\,
            in3 => \N__43828\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6621_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__56065\,
            in1 => \N__44156\,
            in2 => \_gnd_net_\,
            in3 => \N__56451\,
            lcout => n8_adj_1625,
            ltout => \n8_adj_1625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_4_i15_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__63654\,
            in1 => \N__57582\,
            in2 => \N__43798\,
            in3 => \N__44181\,
            lcout => \data_index_9_N_236_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57583\,
            in1 => \N__51339\,
            in2 => \N__46658\,
            in3 => \N__44383\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__47014\,
            in1 => \N__51323\,
            in2 => \N__49133\,
            in3 => \N__57587\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i4_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__44182\,
            in1 => \N__44170\,
            in2 => \N__57701\,
            in3 => \N__63655\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61918\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20577_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__59961\,
            in1 => \N__60478\,
            in2 => \N__56917\,
            in3 => \N__44350\,
            lcout => n23546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_124_Mux_0_i30_4_lut_4_lut_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011110011010"
        )
    port map (
            in0 => \N__60479\,
            in1 => \N__59227\,
            in2 => \N__61018\,
            in3 => \N__59962\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_259_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__49396\,
            in1 => \N__49655\,
            in2 => \N__47013\,
            in3 => \N__49786\,
            lcout => n17_adj_1594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__49656\,
            in1 => \_gnd_net_\,
            in2 => \N__47076\,
            in3 => \N__51363\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48872\,
            in1 => \N__46817\,
            in2 => \_gnd_net_\,
            in3 => \N__44115\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_249_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__44381\,
            in1 => \N__50035\,
            in2 => \N__44079\,
            in3 => \N__50938\,
            lcout => n24_adj_1800,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44078\,
            in1 => \N__51364\,
            in2 => \_gnd_net_\,
            in3 => \N__50808\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20048_2_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44382\,
            lcout => n22314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19242_3_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47391\,
            in1 => \_gnd_net_\,
            in2 => \N__50127\,
            in3 => \N__59009\,
            lcout => n22169,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20387_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__60496\,
            in1 => \N__59536\,
            in2 => \N__46447\,
            in3 => \N__59963\,
            lcout => OPEN,
            ltout => \n23312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23312_bdd_4_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__59965\,
            in1 => \N__44344\,
            in2 => \N__44320\,
            in3 => \N__44288\,
            lcout => OPEN,
            ltout => \n23315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1665080_i1_3_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44188\,
            in2 => \N__44317\,
            in3 => \N__60948\,
            lcout => OPEN,
            ltout => \n30_adj_1741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_3_i127_3_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44314\,
            in2 => \N__44299\,
            in3 => \N__61373\,
            lcout => \comm_buf_1_7_N_559_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57617\,
            in1 => \N__49330\,
            in2 => \N__44295\,
            in3 => \N__46820\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__44272\,
            in1 => \N__59960\,
            in2 => \N__44260\,
            in3 => \N__60495\,
            lcout => OPEN,
            ltout => \n23558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23558_bdd_4_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__44230\,
            in1 => \N__44203\,
            in2 => \N__44191\,
            in3 => \N__59964\,
            lcout => n23561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__44742\,
            in1 => \N__47661\,
            in2 => \N__44764\,
            in3 => \N__44527\,
            lcout => \SIG_DDS.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61971\,
            ce => \N__50404\,
            sr => \N__47674\
        );

    \SIG_DDS.bit_cnt_i2_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__47660\,
            in1 => \_gnd_net_\,
            in2 => \N__44743\,
            in3 => \N__44759\,
            lcout => \SIG_DDS.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61971\,
            ce => \N__50404\,
            sr => \N__47674\
        );

    \SIG_DDS.bit_cnt_i1_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44738\,
            in2 => \_gnd_net_\,
            in3 => \N__47659\,
            lcout => \SIG_DDS.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61971\,
            ce => \N__50404\,
            sr => \N__47674\
        );

    \i16455_2_lut_3_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44715\,
            in1 => \N__62678\,
            in2 => \_gnd_net_\,
            in3 => \N__64076\,
            lcout => n14_adj_1653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16463_2_lut_3_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__64077\,
            in1 => \N__55827\,
            in2 => \N__62690\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16458_2_lut_3_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__64078\,
            in1 => \N__44642\,
            in2 => \N__62691\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__45121\,
            in1 => \N__63742\,
            in2 => \N__57708\,
            in3 => \N__45112\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19893_2_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__44526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50455\,
            lcout => \SIG_DDS.n22671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_9_i15_4_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63738\,
            in1 => \N__44508\,
            in2 => \N__57707\,
            in3 => \N__44496\,
            lcout => \data_index_9_N_236_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6601_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49221\,
            in1 => \N__45135\,
            in2 => \_gnd_net_\,
            in3 => \N__56473\,
            lcout => n8_adj_1621,
            ltout => \n8_adj_1621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_6_i15_4_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57603\,
            in1 => \N__63740\,
            in2 => \N__45115\,
            in3 => \N__45111\,
            lcout => \data_index_9_N_236_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63741\,
            in1 => \N__44926\,
            in2 => \N__57711\,
            in3 => \N__44917\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__44980\,
            in1 => \N__63743\,
            in2 => \N__57709\,
            in3 => \N__44971\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_7_i15_4_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63739\,
            in1 => \N__44925\,
            in2 => \N__57710\,
            in3 => \N__44916\,
            lcout => \data_index_9_N_236_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i0_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000001010101"
        )
    port map (
            in0 => \N__50595\,
            in1 => \N__44812\,
            in2 => \N__44806\,
            in3 => \N__50330\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61996\,
            ce => \N__47632\,
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_16_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50188\,
            in2 => \_gnd_net_\,
            in3 => \N__57119\,
            lcout => \comm_spi.imosi_N_841\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12616_12617_set_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47958\,
            in1 => \N__44783\,
            in2 => \_gnd_net_\,
            in3 => \N__45460\,
            lcout => \comm_spi.n15344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53688\,
            ce => 'H',
            sr => \N__47530\
        );

    \comm_spi.i12604_3_lut_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47954\,
            in1 => \N__44784\,
            in2 => \_gnd_net_\,
            in3 => \N__45458\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i20223_4_lut_3_lut_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45244\,
            in2 => \N__45247\,
            in3 => \N__57070\,
            lcout => \comm_spi.n24019\,
            ltout => \comm_spi.n24019_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12618_3_lut_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__45238\,
            in1 => \N__45232\,
            in2 => \N__45226\,
            in3 => \_gnd_net_\,
            lcout => comm_rx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_112_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47919\,
            in1 => \N__48051\,
            in2 => \N__47833\,
            in3 => \N__48021\,
            lcout => n31_adj_1680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47937\,
            in1 => \N__47868\,
            in2 => \N__47890\,
            in3 => \N__48085\,
            lcout => n33,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_adj_110_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47973\,
            in1 => \N__48235\,
            in2 => \N__48106\,
            in3 => \N__48202\,
            lcout => n32,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_202_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45222\,
            in1 => \N__45208\,
            in2 => \N__45190\,
            in3 => \N__45169\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__60063\,
            in1 => \N__60358\,
            in2 => \_gnd_net_\,
            in3 => \N__59185\,
            lcout => n11379,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47904\,
            in1 => \N__48165\,
            in2 => \N__47854\,
            in3 => \N__48216\,
            lcout => n30_adj_1681,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48135\,
            in1 => \N__48120\,
            in2 => \N__48184\,
            in3 => \N__48150\,
            lcout => OPEN,
            ltout => \n12_adj_1760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48036\,
            in1 => \N__47991\,
            in2 => \N__45496\,
            in3 => \N__48436\,
            lcout => OPEN,
            ltout => \n20834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_109_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__48006\,
            in1 => \N__48066\,
            in2 => \N__45493\,
            in3 => \N__45490\,
            lcout => OPEN,
            ltout => \n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18_4_lut_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45484\,
            in1 => \N__45478\,
            in2 => \N__45472\,
            in3 => \N__45469\,
            lcout => n49,
            ltout => \n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_flag_292_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45463\,
            in3 => \N__52659\,
            lcout => wdtick_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48405\,
            ce => 'H',
            sr => \N__51225\
        );

    \comm_spi.i20208_4_lut_3_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45454\,
            in1 => \N__57049\,
            in2 => \_gnd_net_\,
            in3 => \N__50199\,
            lcout => \comm_spi.n24022\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_66_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46199\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63073\,
            lcout => OPEN,
            ltout => \n8856_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_68_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__57745\,
            in1 => \N__63601\,
            in2 => \N__45430\,
            in3 => \N__59190\,
            lcout => n13273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16182_3_lut_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54527\,
            in1 => \N__55093\,
            in2 => \N__45328\,
            in3 => \_gnd_net_\,
            lcout => n18882,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19916_2_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45727\,
            in2 => \_gnd_net_\,
            in3 => \N__54525\,
            lcout => n22371,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16183_3_lut_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54528\,
            in1 => \_gnd_net_\,
            in2 => \N__45715\,
            in3 => \N__45700\,
            lcout => OPEN,
            ltout => \n18883_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__45667\,
            in1 => \N__45607\,
            in2 => \N__45661\,
            in3 => \N__54307\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61850\,
            ce => \N__46419\,
            sr => \N__46341\
        );

    \i16185_3_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54526\,
            in1 => \N__45625\,
            in2 => \_gnd_net_\,
            in3 => \N__56578\,
            lcout => OPEN,
            ltout => \n18885_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__45616\,
            in1 => \N__54306\,
            in2 => \N__45610\,
            in3 => \N__51800\,
            lcout => n23414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20060_2_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51730\,
            lcout => n22618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i3_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__46257\,
            in1 => \N__62784\,
            in2 => \N__45571\,
            in3 => \N__63595\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_211_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__63594\,
            in1 => \N__45586\,
            in2 => \N__63200\,
            in3 => \N__48301\,
            lcout => n12976,
            ltout => \n12976_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i2_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__54925\,
            in1 => \N__45510\,
            in2 => \N__45520\,
            in3 => \N__63596\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19807_4_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__58950\,
            in1 => \N__60952\,
            in2 => \N__48271\,
            in3 => \N__60396\,
            lcout => OPEN,
            ltout => \n22375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__51514\,
            in1 => \N__63188\,
            in2 => \N__45847\,
            in3 => \N__48642\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_346_Mux_2_i4_3_lut_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__45856\,
            in1 => \N__58210\,
            in2 => \_gnd_net_\,
            in3 => \N__62936\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20075_2_lut_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45844\,
            in2 => \_gnd_net_\,
            in3 => \N__58948\,
            lcout => n22297,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_3787__i3_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__51424\,
            in1 => \N__53771\,
            in2 => \N__51451\,
            in3 => \N__51472\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3787__i3C_net\,
            ce => 'H',
            sr => \N__57122\
        );

    \comm_spi.bit_cnt_3787__i2_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__51471\,
            in1 => \N__51446\,
            in2 => \_gnd_net_\,
            in3 => \N__51423\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3787__i3C_net\,
            ce => 'H',
            sr => \N__57122\
        );

    \comm_spi.bit_cnt_3787__i1_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51470\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3787__i3C_net\,
            ce => 'H',
            sr => \N__57122\
        );

    \comm_spi.bit_cnt_3787__i0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51444\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3787__i3C_net\,
            ce => 'H',
            sr => \N__57122\
        );

    \i12699_2_lut_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45817\,
            in2 => \_gnd_net_\,
            in3 => \N__50020\,
            lcout => n15431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12794_2_lut_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63597\,
            in2 => \_gnd_net_\,
            in3 => \N__45885\,
            lcout => n15517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_226_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46474\,
            in2 => \_gnd_net_\,
            in3 => \N__46520\,
            lcout => n21966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__54792\,
            in1 => \N__46007\,
            in2 => \N__60357\,
            in3 => \N__45949\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16279_2_lut_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60233\,
            in2 => \_gnd_net_\,
            in3 => \N__58840\,
            lcout => n18955,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_332_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__54171\,
            in1 => \N__54068\,
            in2 => \_gnd_net_\,
            in3 => \N__49348\,
            lcout => n12958,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i58_4_lut_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__62530\,
            in1 => \N__45874\,
            in2 => \N__54418\,
            in3 => \N__48901\,
            lcout => n29_adj_1688,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_79_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__58610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50858\,
            lcout => OPEN,
            ltout => \n11402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_133_Mux_2_i127_4_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__55598\,
            in1 => \N__58403\,
            in2 => \N__45859\,
            in3 => \N__61380\,
            lcout => \comm_state_3_N_500_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19773_2_lut_4_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__60902\,
            in1 => \N__58841\,
            in2 => \N__58521\,
            in3 => \N__60247\,
            lcout => n22351,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16149_3_lut_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54542\,
            in1 => \_gnd_net_\,
            in2 => \N__62092\,
            in3 => \N__54949\,
            lcout => OPEN,
            ltout => \n18850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__46210\,
            in1 => \N__46237\,
            in2 => \N__46435\,
            in3 => \N__54331\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61889\,
            ce => \N__46432\,
            sr => \N__46353\
        );

    \i19787_2_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__54539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46276\,
            lcout => n22346,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16150_3_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46258\,
            in1 => \N__46109\,
            in2 => \_gnd_net_\,
            in3 => \N__54541\,
            lcout => n18851,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16152_3_lut_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54540\,
            in1 => \_gnd_net_\,
            in2 => \N__49292\,
            in3 => \N__46228\,
            lcout => OPEN,
            ltout => \n18853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_20444_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__46219\,
            in1 => \N__54330\,
            in2 => \N__46213\,
            in3 => \N__51829\,
            lcout => n23378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16157_3_lut_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__62079\,
            in1 => \N__46200\,
            in2 => \N__46116\,
            in3 => \_gnd_net_\,
            lcout => n18858,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57129\,
            lcout => \comm_spi.data_tx_7__N_874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i7_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46045\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => buf_control_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61905\,
            ce => \N__46687\,
            sr => \N__51646\
        );

    \i1_2_lut_adj_227_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__63050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__64033\,
            lcout => OPEN,
            ltout => \n12021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_291_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__63196\,
            in1 => \N__62675\,
            in2 => \N__46690\,
            in3 => \N__63718\,
            lcout => n12614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i44_3_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__63049\,
            in1 => \N__64031\,
            in2 => \_gnd_net_\,
            in3 => \N__54198\,
            lcout => OPEN,
            ltout => \n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_290_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__63195\,
            in1 => \N__62673\,
            in2 => \N__46681\,
            in3 => \N__63717\,
            lcout => n12548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6984_2_lut_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__62564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63048\,
            lcout => n9714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16459_2_lut_3_lut_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__62674\,
            in1 => \N__46642\,
            in2 => \_gnd_net_\,
            in3 => \N__64032\,
            lcout => n14_adj_1607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_306_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__57712\,
            in1 => \N__46530\,
            in2 => \N__46504\,
            in3 => \N__63650\,
            lcout => n13129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19133_2_lut_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46482\,
            in2 => \_gnd_net_\,
            in3 => \N__58624\,
            lcout => n22059,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_3_i26_3_lut_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__59226\,
            in1 => \_gnd_net_\,
            in2 => \N__47137\,
            in3 => \N__49811\,
            lcout => n26_adj_1740,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_0_i26_3_lut_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47203\,
            in1 => \N__59225\,
            in2 => \_gnd_net_\,
            in3 => \N__49388\,
            lcout => OPEN,
            ltout => \n26_adj_1580_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20582_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__58666\,
            in1 => \N__59974\,
            in2 => \N__47041\,
            in3 => \N__60395\,
            lcout => OPEN,
            ltout => \n23552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23552_bdd_4_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__59975\,
            in1 => \N__47038\,
            in2 => \N__47017\,
            in3 => \N__47009\,
            lcout => n23555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__56022\,
            in1 => \N__51324\,
            in2 => \_gnd_net_\,
            in3 => \N__52481\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61919\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23300_bdd_4_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__46990\,
            in1 => \N__46975\,
            in2 => \N__46960\,
            in3 => \N__59976\,
            lcout => n23303,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19344_3_lut_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46920\,
            in1 => \N__46879\,
            in2 => \_gnd_net_\,
            in3 => \N__60497\,
            lcout => n22271,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19341_3_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59209\,
            in1 => \N__47476\,
            in2 => \_gnd_net_\,
            in3 => \N__49742\,
            lcout => n22268,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__57853\,
            in1 => \N__46851\,
            in2 => \N__52513\,
            in3 => \N__56069\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48879\,
            in1 => \N__46748\,
            in2 => \_gnd_net_\,
            in3 => \N__52625\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i4_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__50769\,
            in1 => \N__57852\,
            in2 => \N__47267\,
            in3 => \N__56070\,
            lcout => buf_dds0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i0_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__57851\,
            in1 => \N__50768\,
            in2 => \N__49140\,
            in3 => \N__47219\,
            lcout => buf_dds0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i0_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__48250\,
            in1 => \N__47202\,
            in2 => \N__63763\,
            in3 => \N__47188\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => n20661,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47175\,
            in1 => \N__52272\,
            in2 => \N__63767\,
            in3 => \N__47161\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n20661,
            carryout => n20662,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47158\,
            in1 => \N__52420\,
            in2 => \N__63764\,
            in3 => \N__47140\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n20662,
            carryout => n20663,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__48942\,
            in1 => \N__47133\,
            in2 => \N__63768\,
            in3 => \N__47119\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n20663,
            carryout => n20664,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__56023\,
            in1 => \N__52563\,
            in2 => \N__63765\,
            in3 => \N__47116\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n20664,
            carryout => n20665,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47099\,
            in1 => \N__51999\,
            in2 => \N__63769\,
            in3 => \N__47080\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n20665,
            carryout => n20666,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47069\,
            in1 => \N__49605\,
            in2 => \N__63766\,
            in3 => \N__47044\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n20666,
            carryout => n20667,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47516\,
            in1 => \N__54672\,
            in2 => \N__63770\,
            in3 => \N__47479\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n20667,
            carryout => n20668,
            clk => \N__61955\,
            ce => \N__47692\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__48871\,
            in1 => \N__47475\,
            in2 => \N__63779\,
            in3 => \N__47461\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => n20669,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__50797\,
            in1 => \N__63748\,
            in2 => \N__50953\,
            in3 => \N__47458\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n20669,
            carryout => n20670,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47451\,
            in1 => \N__47392\,
            in2 => \N__63780\,
            in3 => \N__47380\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n20670,
            carryout => n20671,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__56834\,
            in1 => \N__63752\,
            in2 => \N__56157\,
            in3 => \N__47377\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n20671,
            carryout => n20672,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47352\,
            in1 => \N__49719\,
            in2 => \N__63781\,
            in3 => \N__47317\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n20672,
            carryout => n20673,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__55287\,
            in1 => \N__63756\,
            in2 => \N__61095\,
            in3 => \N__47314\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n20673,
            carryout => n20674,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__51501\,
            in1 => \N__49026\,
            in2 => \N__63782\,
            in3 => \N__47311\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n20674,
            carryout => n20675,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47308\,
            in1 => \N__63760\,
            in2 => \N__47289\,
            in3 => \N__47296\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61972\,
            ce => \N__47691\,
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__52587\,
            in1 => \N__63761\,
            in2 => \N__57855\,
            in3 => \N__53152\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61985\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i20157_4_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__50610\,
            in1 => \N__50536\,
            in2 => \N__47582\,
            in3 => \N__50314\,
            lcout => \SIG_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110111"
        )
    port map (
            in0 => \N__63744\,
            in1 => \N__56479\,
            in2 => \N__57854\,
            in3 => \N__47788\,
            lcout => n13052,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i12835_3_lut_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__50609\,
            in1 => \N__50535\,
            in2 => \_gnd_net_\,
            in3 => \N__50315\,
            lcout => n15562,
            ltout => \n15562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i0_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__50316\,
            in1 => \_gnd_net_\,
            in2 => \N__47665\,
            in3 => \N__47655\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61985\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i1_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50537\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61997\,
            ce => \N__47625\,
            sr => \N__50405\
        );

    \SIG_DDS.SCLK_27_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001010110001"
        )
    port map (
            in0 => \N__50594\,
            in1 => \N__50491\,
            in2 => \N__47601\,
            in3 => \N__50318\,
            lcout => \DDS_SCK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i23_4_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011011"
        )
    port map (
            in0 => \N__50593\,
            in1 => \N__50490\,
            in2 => \N__47583\,
            in3 => \N__50317\,
            lcout => \SIG_DDS.n9_adj_1490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_17_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57096\,
            lcout => \comm_spi.DOUT_7__N_834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12602_12603_set_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50198\,
            lcout => \comm_spi.n15330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61832\,
            ce => 'H',
            sr => \N__50140\
        );

    \wdtick_cnt_3783_3784__i1_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48541\,
            in1 => \N__47938\,
            in2 => \_gnd_net_\,
            in3 => \N__47923\,
            lcout => wdtick_cnt_0,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => n20766,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48510\,
            in1 => \N__47920\,
            in2 => \_gnd_net_\,
            in3 => \N__47908\,
            lcout => wdtick_cnt_1,
            ltout => OPEN,
            carryin => n20766,
            carryout => n20767,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i3_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48542\,
            in1 => \N__47905\,
            in2 => \_gnd_net_\,
            in3 => \N__47893\,
            lcout => wdtick_cnt_2,
            ltout => OPEN,
            carryin => n20767,
            carryout => n20768,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i4_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48511\,
            in1 => \N__47883\,
            in2 => \_gnd_net_\,
            in3 => \N__47872\,
            lcout => wdtick_cnt_3,
            ltout => OPEN,
            carryin => n20768,
            carryout => n20769,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i5_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48543\,
            in1 => \N__47869\,
            in2 => \_gnd_net_\,
            in3 => \N__47857\,
            lcout => wdtick_cnt_4,
            ltout => OPEN,
            carryin => n20769,
            carryout => n20770,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i6_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48512\,
            in1 => \N__47847\,
            in2 => \_gnd_net_\,
            in3 => \N__47836\,
            lcout => wdtick_cnt_5,
            ltout => OPEN,
            carryin => n20770,
            carryout => n20771,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i7_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48544\,
            in1 => \N__47832\,
            in2 => \_gnd_net_\,
            in3 => \N__47818\,
            lcout => wdtick_cnt_6,
            ltout => OPEN,
            carryin => n20771,
            carryout => n20772,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i8_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48513\,
            in1 => \N__48099\,
            in2 => \_gnd_net_\,
            in3 => \N__48088\,
            lcout => wdtick_cnt_7,
            ltout => OPEN,
            carryin => n20772,
            carryout => n20773,
            clk => \N__48406\,
            ce => \N__48349\,
            sr => \N__51226\
        );

    \wdtick_cnt_3783_3784__i9_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48505\,
            in1 => \N__48084\,
            in2 => \_gnd_net_\,
            in3 => \N__48070\,
            lcout => wdtick_cnt_8,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => n20774,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i10_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48533\,
            in1 => \N__48067\,
            in2 => \_gnd_net_\,
            in3 => \N__48055\,
            lcout => wdtick_cnt_9,
            ltout => OPEN,
            carryin => n20774,
            carryout => n20775,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i11_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48502\,
            in1 => \N__48052\,
            in2 => \_gnd_net_\,
            in3 => \N__48040\,
            lcout => wdtick_cnt_10,
            ltout => OPEN,
            carryin => n20775,
            carryout => n20776,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i12_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48534\,
            in1 => \N__48037\,
            in2 => \_gnd_net_\,
            in3 => \N__48025\,
            lcout => wdtick_cnt_11,
            ltout => OPEN,
            carryin => n20776,
            carryout => n20777,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i13_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48503\,
            in1 => \N__48022\,
            in2 => \_gnd_net_\,
            in3 => \N__48010\,
            lcout => wdtick_cnt_12,
            ltout => OPEN,
            carryin => n20777,
            carryout => n20778,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i14_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48535\,
            in1 => \N__48007\,
            in2 => \_gnd_net_\,
            in3 => \N__47995\,
            lcout => wdtick_cnt_13,
            ltout => OPEN,
            carryin => n20778,
            carryout => n20779,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i15_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48504\,
            in1 => \N__47992\,
            in2 => \_gnd_net_\,
            in3 => \N__47977\,
            lcout => wdtick_cnt_14,
            ltout => OPEN,
            carryin => n20779,
            carryout => n20780,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i16_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48536\,
            in1 => \N__47974\,
            in2 => \_gnd_net_\,
            in3 => \N__47962\,
            lcout => wdtick_cnt_15,
            ltout => OPEN,
            carryin => n20780,
            carryout => n20781,
            clk => \N__48407\,
            ce => \N__48338\,
            sr => \N__51224\
        );

    \wdtick_cnt_3783_3784__i17_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48537\,
            in1 => \N__48234\,
            in2 => \_gnd_net_\,
            in3 => \N__48220\,
            lcout => wdtick_cnt_16,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => n20782,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i18_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48506\,
            in1 => \N__48217\,
            in2 => \_gnd_net_\,
            in3 => \N__48205\,
            lcout => wdtick_cnt_17,
            ltout => OPEN,
            carryin => n20782,
            carryout => n20783,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i19_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48538\,
            in1 => \N__48201\,
            in2 => \_gnd_net_\,
            in3 => \N__48187\,
            lcout => wdtick_cnt_18,
            ltout => OPEN,
            carryin => n20783,
            carryout => n20784,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i20_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48507\,
            in1 => \N__48183\,
            in2 => \_gnd_net_\,
            in3 => \N__48169\,
            lcout => wdtick_cnt_19,
            ltout => OPEN,
            carryin => n20784,
            carryout => n20785,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i21_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48539\,
            in1 => \N__48166\,
            in2 => \_gnd_net_\,
            in3 => \N__48154\,
            lcout => wdtick_cnt_20,
            ltout => OPEN,
            carryin => n20785,
            carryout => n20786,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i22_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48508\,
            in1 => \N__48151\,
            in2 => \_gnd_net_\,
            in3 => \N__48139\,
            lcout => wdtick_cnt_21,
            ltout => OPEN,
            carryin => n20786,
            carryout => n20787,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i23_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48540\,
            in1 => \N__48136\,
            in2 => \_gnd_net_\,
            in3 => \N__48124\,
            lcout => wdtick_cnt_22,
            ltout => OPEN,
            carryin => n20787,
            carryout => n20788,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i24_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__48509\,
            in1 => \N__48121\,
            in2 => \_gnd_net_\,
            in3 => \N__48109\,
            lcout => wdtick_cnt_23,
            ltout => OPEN,
            carryin => n20788,
            carryout => n20789,
            clk => \N__48408\,
            ce => \N__48337\,
            sr => \N__51219\
        );

    \wdtick_cnt_3783_3784__i25_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__48435\,
            in1 => \N__48532\,
            in2 => \_gnd_net_\,
            in3 => \N__48439\,
            lcout => wdtick_cnt_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48410\,
            ce => \N__48345\,
            sr => \N__51223\
        );

    \i2_2_lut_4_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__51168\,
            in1 => \N__51784\,
            in2 => \N__62608\,
            in3 => \N__57353\,
            lcout => n7_adj_1757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__58042\,
            in1 => \N__58208\,
            in2 => \N__51808\,
            in3 => \N__54310\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61865\,
            ce => \N__48262\,
            sr => \N__48292\
        );

    \i462_2_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58040\,
            lcout => n2562,
            ltout => \n2562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i2_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__51785\,
            in1 => \N__54309\,
            in2 => \N__48295\,
            in3 => \N__54572\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61865\,
            ce => \N__48262\,
            sr => \N__48292\
        );

    \comm_index_i0_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__58207\,
            in1 => \N__54308\,
            in2 => \_gnd_net_\,
            in3 => \N__58041\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61865\,
            ce => \N__48262\,
            sr => \N__48292\
        );

    \i3_3_lut_4_lut_adj_284_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__61381\,
            in1 => \N__60006\,
            in2 => \N__64066\,
            in3 => \N__63505\,
            lcout => n8_adj_1782,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_286_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__63504\,
            in1 => \N__51175\,
            in2 => \_gnd_net_\,
            in3 => \N__63204\,
            lcout => n12540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_78_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__64034\,
            in1 => \N__49087\,
            in2 => \_gnd_net_\,
            in3 => \N__62449\,
            lcout => n14_adj_1606,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19313_4_lut_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__64023\,
            in1 => \N__53439\,
            in2 => \N__48673\,
            in3 => \N__48655\,
            lcout => OPEN,
            ltout => \n22240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57739\,
            in2 => \N__48658\,
            in3 => \N__63494\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61878\,
            ce => \N__51235\,
            sr => \_gnd_net_\
        );

    \i20126_3_lut_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__62572\,
            in1 => \N__57300\,
            in2 => \_gnd_net_\,
            in3 => \N__51169\,
            lcout => n23053,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12533_2_lut_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58153\,
            in2 => \_gnd_net_\,
            in3 => \N__62930\,
            lcout => n15261,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_128_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__62931\,
            in1 => \N__62570\,
            in2 => \_gnd_net_\,
            in3 => \N__64022\,
            lcout => OPEN,
            ltout => \n11280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_228_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__63492\,
            in1 => \N__63145\,
            in2 => \N__48649\,
            in3 => \N__56247\,
            lcout => n12509,
            ltout => \n12509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_114_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__64024\,
            in1 => \N__62571\,
            in2 => \N__48646\,
            in3 => \N__63493\,
            lcout => n18363,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_86_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__54312\,
            in1 => \N__48643\,
            in2 => \N__48628\,
            in3 => \N__54537\,
            lcout => n4_adj_1745,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23486_bdd_4_lut_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__48609\,
            in1 => \N__48586\,
            in2 => \N__48574\,
            in3 => \N__60309\,
            lcout => n22180,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_311_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51133\,
            in3 => \N__54538\,
            lcout => n4_adj_1749,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19973_2_lut_4_lut_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110111"
        )
    port map (
            in0 => \N__58650\,
            in1 => \N__60314\,
            in2 => \N__50885\,
            in3 => \N__59015\,
            lcout => n22330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i50_4_lut_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101101010000"
        )
    port map (
            in0 => \N__59014\,
            in1 => \N__59867\,
            in2 => \N__60463\,
            in3 => \N__60990\,
            lcout => OPEN,
            ltout => \n46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19794_4_lut_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__58649\,
            in1 => \N__59887\,
            in2 => \N__48997\,
            in3 => \N__60313\,
            lcout => n22353,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_0_i111_3_lut_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__59016\,
            in1 => \_gnd_net_\,
            in2 => \N__48994\,
            in3 => \N__48964\,
            lcout => n111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_323_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__62905\,
            in1 => \N__54311\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16444_2_lut_3_lut_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__62567\,
            in1 => \N__49273\,
            in2 => \_gnd_net_\,
            in3 => \N__64030\,
            lcout => n14_adj_1662,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_312_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100010001"
        )
    port map (
            in0 => \N__51623\,
            in1 => \N__62565\,
            in2 => \N__49362\,
            in3 => \N__48900\,
            lcout => n12_adj_1684,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i0_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48880\,
            in1 => \N__48798\,
            in2 => \_gnd_net_\,
            in3 => \N__48692\,
            lcout => \buf_cfgRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16282_2_lut_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58515\,
            in2 => \_gnd_net_\,
            in3 => \N__58625\,
            lcout => n7148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_297_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__58626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59936\,
            lcout => OPEN,
            ltout => \n4_adj_1709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i45_4_lut_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__49372\,
            in1 => \N__58399\,
            in2 => \N__49366\,
            in3 => \N__61379\,
            lcout => n30_adj_1720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19163_2_lut_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__54326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62943\,
            lcout => n22089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_330_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100010001"
        )
    port map (
            in0 => \N__51624\,
            in1 => \N__62566\,
            in2 => \N__49363\,
            in3 => \N__51585\,
            lcout => n12_adj_1802,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62598\,
            in1 => \N__62788\,
            in2 => \_gnd_net_\,
            in3 => \N__49342\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61920\,
            ce => \N__55769\,
            sr => \N__55707\
        );

    \comm_buf_1__i6_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__53883\,
            in1 => \N__62599\,
            in2 => \_gnd_net_\,
            in3 => \N__49615\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61920\,
            ce => \N__55769\,
            sr => \N__55707\
        );

    \comm_buf_1__i0_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62597\,
            in1 => \N__54023\,
            in2 => \_gnd_net_\,
            in3 => \N__51655\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61920\,
            ce => \N__55769\,
            sr => \N__55707\
        );

    \i19785_2_lut_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49030\,
            in2 => \_gnd_net_\,
            in3 => \N__59191\,
            lcout => n22296,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19894_2_lut_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__59192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49723\,
            lcout => n22499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23516_bdd_4_lut_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__49690\,
            in1 => \N__59978\,
            in2 => \N__49669\,
            in3 => \N__49588\,
            lcout => OPEN,
            ltout => \n23519_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1668899_i1_3_lut_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60976\,
            in1 => \_gnd_net_\,
            in2 => \N__49642\,
            in3 => \N__49639\,
            lcout => OPEN,
            ltout => \n30_adj_1724_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_6_i127_3_lut_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49627\,
            in2 => \N__49618\,
            in3 => \N__61383\,
            lcout => \comm_buf_1_7_N_559_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_6_i26_3_lut_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49609\,
            in1 => \N__59502\,
            in2 => \_gnd_net_\,
            in3 => \N__49778\,
            lcout => OPEN,
            ltout => \n26_adj_1723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20572_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__55441\,
            in1 => \N__59977\,
            in2 => \N__49591\,
            in3 => \N__60603\,
            lcout => n23516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16700105_i1_3_lut_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60975\,
            in1 => \N__49582\,
            in2 => \_gnd_net_\,
            in3 => \N__49576\,
            lcout => n30_adj_1579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i4_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__49457\,
            in1 => \N__55381\,
            in2 => \N__56086\,
            in3 => \N__49502\,
            lcout => buf_dds1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49392\,
            in2 => \N__49438\,
            in3 => \_gnd_net_\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => n20622,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i1_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52257\,
            in2 => \_gnd_net_\,
            in3 => \N__49825\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n20622,
            carryout => n20623,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i2_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52398\,
            in2 => \_gnd_net_\,
            in3 => \N__49822\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n20623,
            carryout => n20624,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i3_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49815\,
            in2 => \_gnd_net_\,
            in3 => \N__49795\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n20624,
            carryout => n20625,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i4_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52545\,
            in2 => \_gnd_net_\,
            in3 => \N__49792\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n20625,
            carryout => n20626,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i5_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51980\,
            in2 => \_gnd_net_\,
            in3 => \N__49789\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n20626,
            carryout => n20627,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i6_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49782\,
            in2 => \_gnd_net_\,
            in3 => \N__49762\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n20627,
            carryout => n20628,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i7_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54650\,
            in2 => \_gnd_net_\,
            in3 => \N__49759\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n20628,
            carryout => n20629,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__50018\,
            sr => \N__49942\
        );

    \data_cntvec_i0_i8_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49746\,
            in2 => \_gnd_net_\,
            in3 => \N__49726\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => n20630,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i9_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50937\,
            in2 => \_gnd_net_\,
            in3 => \N__50131\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n20630,
            carryout => n20631,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i10_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50117\,
            in2 => \_gnd_net_\,
            in3 => \N__50092\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n20631,
            carryout => n20632,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i11_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56132\,
            in2 => \_gnd_net_\,
            in3 => \N__50089\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n20632,
            carryout => n20633,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i12_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50082\,
            in2 => \_gnd_net_\,
            in3 => \N__50068\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n20633,
            carryout => n20634,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i13_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50058\,
            in2 => \_gnd_net_\,
            in3 => \N__50044\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n20634,
            carryout => n20635,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i14_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51699\,
            in2 => \_gnd_net_\,
            in3 => \N__50041\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n20635,
            carryout => n20636,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \data_cntvec_i0_i15_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50034\,
            in2 => \_gnd_net_\,
            in3 => \N__50038\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__50017\,
            sr => \N__49943\
        );

    \n23480_bdd_4_lut_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__49909\,
            in1 => \N__60592\,
            in2 => \N__49884\,
            in3 => \N__49852\,
            lcout => OPEN,
            ltout => \n22183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_20528_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__61022\,
            in1 => \N__60059\,
            in2 => \N__49828\,
            in3 => \N__50899\,
            lcout => OPEN,
            ltout => \n23462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23462_bdd_4_lut_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__50986\,
            in1 => \N__50977\,
            in2 => \N__50968\,
            in3 => \N__61023\,
            lcout => n23465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19257_3_lut_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50949\,
            in1 => \N__59408\,
            in2 => \_gnd_net_\,
            in3 => \N__50933\,
            lcout => OPEN,
            ltout => \n22184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19259_4_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__59409\,
            in1 => \N__50917\,
            in2 => \N__50902\,
            in3 => \N__60591\,
            lcout => n22186,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_285_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__60058\,
            in1 => \N__58528\,
            in2 => \_gnd_net_\,
            in3 => \N__61021\,
            lcout => n21997,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i9_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50807\,
            in1 => \N__50633\,
            in2 => \_gnd_net_\,
            in3 => \N__50775\,
            lcout => buf_dds0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.CS_28_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__50608\,
            in1 => \N__50538\,
            in2 => \_gnd_net_\,
            in3 => \N__50329\,
            lcout => \DDS_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__62008\,
            ce => \N__50245\,
            sr => \_gnd_net_\
        );

    \i20042_2_lut_LC_18_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50233\,
            in2 => \_gnd_net_\,
            in3 => \N__59427\,
            lcout => n22595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_18_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57077\,
            lcout => \comm_spi.imosi_N_840\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12628_12629_reset_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51124\,
            in1 => \N__51103\,
            in2 => \_gnd_net_\,
            in3 => \N__51079\,
            lcout => \comm_spi.n15357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53670\,
            ce => 'H',
            sr => \N__51022\
        );

    \i19790_2_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56871\,
            in2 => \_gnd_net_\,
            in3 => \N__63030\,
            lcout => OPEN,
            ltout => \n22489_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001110101"
        )
    port map (
            in0 => \N__63358\,
            in1 => \N__57521\,
            in2 => \N__51004\,
            in3 => \N__50992\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61866\,
            ce => \N__50998\,
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__62485\,
            in1 => \N__63029\,
            in2 => \N__54183\,
            in3 => \N__57354\,
            lcout => OPEN,
            ltout => \n20959_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_88_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__57970\,
            in1 => \N__51566\,
            in2 => \N__51001\,
            in3 => \N__53349\,
            lcout => n21883,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_70_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64006\,
            in2 => \_gnd_net_\,
            in3 => \N__63357\,
            lcout => n12951,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_346_Mux_3_i7_4_lut_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__62486\,
            in1 => \N__51406\,
            in2 => \N__53416\,
            in3 => \N__64007\,
            lcout => n19241,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19824_2_lut_3_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__58117\,
            in1 => \N__62421\,
            in2 => \_gnd_net_\,
            in3 => \N__58036\,
            lcout => n22339,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111101111"
        )
    port map (
            in0 => \N__58037\,
            in1 => \N__58118\,
            in2 => \N__62601\,
            in3 => \N__62933\,
            lcout => n22033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_304_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__53438\,
            in1 => \N__62427\,
            in2 => \N__54184\,
            in3 => \N__58038\,
            lcout => OPEN,
            ltout => \n12064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_143_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__51244\,
            in1 => \N__51567\,
            in2 => \N__51238\,
            in3 => \N__53350\,
            lcout => n21885,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19147_2_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__62934\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62426\,
            lcout => OPEN,
            ltout => \n22073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_224_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000100"
        )
    port map (
            in0 => \N__64011\,
            in1 => \N__63173\,
            in2 => \N__51229\,
            in3 => \N__63378\,
            lcout => n12050,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \flagcntwd_306_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__62935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62428\,
            lcout => flagcntwd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61879\,
            ce => \N__51184\,
            sr => \N__51645\
        );

    \i17_3_lut_3_lut_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__62422\,
            in1 => \_gnd_net_\,
            in2 => \N__64050\,
            in3 => \N__62932\,
            lcout => n10_adj_1602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_106_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__51780\,
            in1 => \N__51166\,
            in2 => \N__58181\,
            in3 => \N__58018\,
            lcout => n21956,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_107_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__51167\,
            in1 => \N__58151\,
            in2 => \N__58039\,
            in3 => \N__51779\,
            lcout => n29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12123_2_lut_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__62569\,
            in1 => \N__62906\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n14851,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__58152\,
            in1 => \N__62568\,
            in2 => \_gnd_net_\,
            in3 => \N__51568\,
            lcout => n21981,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_132_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__53398\,
            in1 => \N__63985\,
            in2 => \N__51547\,
            in3 => \N__63613\,
            lcout => n11_adj_1585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__51502\,
            in1 => \N__51283\,
            in2 => \N__51729\,
            in3 => \_gnd_net_\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__51469\,
            in1 => \N__51450\,
            in2 => \_gnd_net_\,
            in3 => \N__51422\,
            lcout => \comm_spi.n18536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19781_2_lut_3_lut_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__62907\,
            in1 => \N__58147\,
            in2 => \_gnd_net_\,
            in3 => \N__57299\,
            lcout => n22487,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_52_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__63393\,
            in1 => \N__51397\,
            in2 => \N__57763\,
            in3 => \N__58369\,
            lcout => n13171,
            ltout => \n13171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57953\,
            in2 => \N__51247\,
            in3 => \N__56838\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20051_2_lut_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58526\,
            in2 => \_gnd_net_\,
            in3 => \N__58651\,
            lcout => n22329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_326_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__54445\,
            in3 => \N__54546\,
            lcout => n20318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_130_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__51877\,
            in1 => \N__58527\,
            in2 => \N__51865\,
            in3 => \N__61362\,
            lcout => \comm_state_3_N_484_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_87_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__51856\,
            in1 => \N__51844\,
            in2 => \_gnd_net_\,
            in3 => \N__51807\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_251_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__51725\,
            in1 => \N__51703\,
            in2 => \N__57957\,
            in3 => \N__56137\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11570_3_lut_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__61363\,
            in1 => \N__51670\,
            in2 => \_gnd_net_\,
            in3 => \N__51664\,
            lcout => \comm_buf_1_7_N_559_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_82_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__62481\,
            in1 => \N__63994\,
            in2 => \_gnd_net_\,
            in3 => \N__63382\,
            lcout => n21271,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_317_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__62596\,
            in1 => \N__51625\,
            in2 => \N__51601\,
            in3 => \N__51589\,
            lcout => OPEN,
            ltout => \n12_adj_1677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_318_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__54160\,
            in1 => \_gnd_net_\,
            in2 => \N__51574\,
            in3 => \N__54066\,
            lcout => n12892,
            ltout => \n12892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12787_2_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__63381\,
            in1 => \_gnd_net_\,
            in2 => \N__51571\,
            in3 => \_gnd_net_\,
            lcout => n15510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_209_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__62480\,
            in1 => \N__63993\,
            in2 => \_gnd_net_\,
            in3 => \N__63379\,
            lcout => n12966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i72_4_lut_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__62595\,
            in1 => \N__58378\,
            in2 => \N__54417\,
            in3 => \N__54430\,
            lcout => OPEN,
            ltout => \n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_301_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__54159\,
            in1 => \N__54067\,
            in2 => \N__52009\,
            in3 => \N__62969\,
            lcout => n12761,
            ltout => \n12761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12766_2_lut_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__63380\,
            in1 => \_gnd_net_\,
            in2 => \N__52006\,
            in3 => \_gnd_net_\,
            lcout => n15489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_5_i26_3_lut_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59505\,
            in1 => \N__52003\,
            in2 => \_gnd_net_\,
            in3 => \N__51981\,
            lcout => OPEN,
            ltout => \n26_adj_1730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20414_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__59554\,
            in1 => \N__59982\,
            in2 => \N__51958\,
            in3 => \N__60521\,
            lcout => OPEN,
            ltout => \n23336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23336_bdd_4_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__59984\,
            in1 => \N__51955\,
            in2 => \N__51928\,
            in3 => \N__51924\,
            lcout => OPEN,
            ltout => \n23339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1668296_i1_3_lut_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52282\,
            in2 => \N__51901\,
            in3 => \N__60957\,
            lcout => OPEN,
            ltout => \n30_adj_1731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_5_i127_3_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61408\,
            in2 => \N__51898\,
            in3 => \N__51895\,
            lcout => OPEN,
            ltout => \comm_buf_1_7_N_559_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__55170\,
            in1 => \N__62600\,
            in2 => \N__52363\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61941\,
            ce => \N__55751\,
            sr => \N__55714\
        );

    \n23354_bdd_4_lut_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__59983\,
            in1 => \N__52360\,
            in2 => \N__52342\,
            in3 => \N__52297\,
            lcout => n23357,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_1_i26_3_lut_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__52276\,
            in1 => \N__59503\,
            in2 => \_gnd_net_\,
            in3 => \N__52247\,
            lcout => n26_adj_1753,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19215_3_lut_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60519\,
            in1 => \N__52234\,
            in2 => \_gnd_net_\,
            in3 => \N__52207\,
            lcout => OPEN,
            ltout => \n22142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_20468_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__60977\,
            in1 => \N__59987\,
            in2 => \N__52183\,
            in3 => \N__52015\,
            lcout => OPEN,
            ltout => \n23408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23408_bdd_4_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__52180\,
            in1 => \N__52681\,
            in2 => \N__52162\,
            in3 => \N__60978\,
            lcout => OPEN,
            ltout => \n23411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_1_i127_3_lut_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61407\,
            in2 => \N__52159\,
            in3 => \N__52156\,
            lcout => OPEN,
            ltout => \comm_buf_1_7_N_559_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i1_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__54796\,
            in1 => \_gnd_net_\,
            in2 => \N__52147\,
            in3 => \N__62671\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61957\,
            ce => \N__55767\,
            sr => \N__55709\
        );

    \i19216_4_lut_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__52039\,
            in1 => \N__60518\,
            in2 => \N__52024\,
            in3 => \N__59504\,
            lcout => n22143,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_4_i26_3_lut_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__52567\,
            in1 => \N__59506\,
            in2 => \_gnd_net_\,
            in3 => \N__52541\,
            lcout => OPEN,
            ltout => \n26_adj_1735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20400_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__52525\,
            in1 => \N__59985\,
            in2 => \N__52516\,
            in3 => \N__60520\,
            lcout => OPEN,
            ltout => \n23318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23318_bdd_4_lut_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__59986\,
            in1 => \N__52512\,
            in2 => \N__52489\,
            in3 => \N__52486\,
            lcout => OPEN,
            ltout => \n23321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1667693_i1_3_lut_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52462\,
            in2 => \N__52447\,
            in3 => \N__60979\,
            lcout => OPEN,
            ltout => \n30_adj_1736_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_4_i127_3_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52444\,
            in2 => \N__52426\,
            in3 => \N__61352\,
            lcout => OPEN,
            ltout => \comm_buf_1_7_N_559_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__55060\,
            in1 => \_gnd_net_\,
            in2 => \N__52423\,
            in3 => \N__62670\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61974\,
            ce => \N__55768\,
            sr => \N__55700\
        );

    \mux_126_Mux_2_i26_3_lut_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__52419\,
            in1 => \N__59507\,
            in2 => \_gnd_net_\,
            in3 => \N__52397\,
            lcout => OPEN,
            ltout => \n26_adj_1748_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19225_4_lut_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__59508\,
            in1 => \N__52378\,
            in2 => \N__52366\,
            in3 => \N__60647\,
            lcout => OPEN,
            ltout => \n22152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_20493_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__52786\,
            in1 => \N__60065\,
            in2 => \N__52993\,
            in3 => \N__61024\,
            lcout => OPEN,
            ltout => \n23444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23444_bdd_4_lut_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__61025\,
            in1 => \N__52990\,
            in2 => \N__52972\,
            in3 => \N__52969\,
            lcout => OPEN,
            ltout => \n23447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_2_i127_3_lut_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52957\,
            in2 => \N__52942\,
            in3 => \N__61411\,
            lcout => OPEN,
            ltout => \comm_buf_1_7_N_559_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54929\,
            in2 => \N__52939\,
            in3 => \N__62672\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61986\,
            ce => \N__55774\,
            sr => \N__55708\
        );

    \i19224_3_lut_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__60646\,
            in1 => \N__52843\,
            in2 => \_gnd_net_\,
            in3 => \N__52812\,
            lcout => n22151,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i23_3_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__52779\,
            in1 => \N__59410\,
            in2 => \_gnd_net_\,
            in3 => \N__52744\,
            lcout => n23_adj_1791,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19209_3_lut_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52716\,
            in1 => \N__52690\,
            in2 => \_gnd_net_\,
            in3 => \N__60593\,
            lcout => n22136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16252_2_lut_2_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52669\,
            in2 => \_gnd_net_\,
            in3 => \N__52638\,
            lcout => \CONT_SD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_0_i15_4_lut_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__63525\,
            in1 => \N__52588\,
            in2 => \N__57872\,
            in3 => \N__53151\,
            lcout => \data_index_9_N_236_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20091_2_lut_LC_19_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53035\,
            in2 => \_gnd_net_\,
            in3 => \N__59399\,
            lcout => n22500,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0on_i0_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56722\,
            in2 => \_gnd_net_\,
            in3 => \N__53014\,
            lcout => \ADC_VDC.genclk.t0on_0\,
            ltout => OPEN,
            carryin => \bfn_19_5_0_\,
            carryout => \ADC_VDC.genclk.n20751\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i1_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56752\,
            in2 => \N__64844\,
            in3 => \N__53011\,
            lcout => \ADC_VDC.genclk.t0on_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20751\,
            carryout => \ADC_VDC.genclk.n20752\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i2_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64780\,
            in2 => \N__56692\,
            in3 => \N__53008\,
            lcout => \ADC_VDC.genclk.t0on_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20752\,
            carryout => \ADC_VDC.genclk.n20753\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i3_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57244\,
            in2 => \N__64845\,
            in3 => \N__53005\,
            lcout => \ADC_VDC.genclk.t0on_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20753\,
            carryout => \ADC_VDC.genclk.n20754\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i4_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64784\,
            in2 => \N__56740\,
            in3 => \N__53002\,
            lcout => \ADC_VDC.genclk.t0on_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20754\,
            carryout => \ADC_VDC.genclk.n20755\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i5_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57231\,
            in2 => \N__64846\,
            in3 => \N__52999\,
            lcout => \ADC_VDC.genclk.t0on_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20755\,
            carryout => \ADC_VDC.genclk.n20756\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i6_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64788\,
            in2 => \N__56767\,
            in3 => \N__52996\,
            lcout => \ADC_VDC.genclk.t0on_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20756\,
            carryout => \ADC_VDC.genclk.n20757\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i7_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56676\,
            in2 => \N__64847\,
            in3 => \N__53179\,
            lcout => \ADC_VDC.genclk.t0on_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20757\,
            carryout => \ADC_VDC.genclk.n20758\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57199\,
            sr => \N__64447\
        );

    \ADC_VDC.genclk.t0on_i8_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57217\,
            in2 => \N__64696\,
            in3 => \N__53176\,
            lcout => \ADC_VDC.genclk.t0on_8\,
            ltout => OPEN,
            carryin => \bfn_19_6_0_\,
            carryout => \ADC_VDC.genclk.n20759\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i9_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64641\,
            in2 => \N__56632\,
            in3 => \N__53173\,
            lcout => \ADC_VDC.genclk.t0on_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20759\,
            carryout => \ADC_VDC.genclk.n20760\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i10_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56662\,
            in2 => \N__64693\,
            in3 => \N__53170\,
            lcout => \ADC_VDC.genclk.t0on_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20760\,
            carryout => \ADC_VDC.genclk.n20761\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i11_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64629\,
            in2 => \N__56602\,
            in3 => \N__53167\,
            lcout => \ADC_VDC.genclk.t0on_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20761\,
            carryout => \ADC_VDC.genclk.n20762\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i12_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56706\,
            in2 => \N__64694\,
            in3 => \N__53164\,
            lcout => \ADC_VDC.genclk.t0on_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20762\,
            carryout => \ADC_VDC.genclk.n20763\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i13_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64633\,
            in2 => \N__57262\,
            in3 => \N__53161\,
            lcout => \ADC_VDC.genclk.t0on_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20763\,
            carryout => \ADC_VDC.genclk.n20764\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i14_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56644\,
            in2 => \N__64695\,
            in3 => \N__53158\,
            lcout => \ADC_VDC.genclk.t0on_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20764\,
            carryout => \ADC_VDC.genclk.n20765\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \ADC_VDC.genclk.t0on_i15_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56616\,
            in1 => \N__64637\,
            in2 => \_gnd_net_\,
            in3 => \N__53155\,
            lcout => \ADC_VDC.genclk.t0on_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57195\,
            sr => \N__64457\
        );

    \dds0_mclkcnt_i7_3792__i0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53245\,
            in2 => \_gnd_net_\,
            in3 => \N__53209\,
            lcout => dds0_mclkcnt_0,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => n20819,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53286\,
            in2 => \_gnd_net_\,
            in3 => \N__53206\,
            lcout => dds0_mclkcnt_1,
            ltout => OPEN,
            carryin => n20819,
            carryout => n20820,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53230\,
            in2 => \_gnd_net_\,
            in3 => \N__53203\,
            lcout => dds0_mclkcnt_2,
            ltout => OPEN,
            carryin => n20820,
            carryout => n20821,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53314\,
            in2 => \_gnd_net_\,
            in3 => \N__53200\,
            lcout => dds0_mclkcnt_3,
            ltout => OPEN,
            carryin => n20821,
            carryout => n20822,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53272\,
            in2 => \_gnd_net_\,
            in3 => \N__53197\,
            lcout => dds0_mclkcnt_4,
            ltout => OPEN,
            carryin => n20822,
            carryout => n20823,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53302\,
            in2 => \_gnd_net_\,
            in3 => \N__53194\,
            lcout => dds0_mclkcnt_5,
            ltout => OPEN,
            carryin => n20823,
            carryout => n20824,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53185\,
            in2 => \_gnd_net_\,
            in3 => \N__53191\,
            lcout => dds0_mclkcnt_6,
            ltout => OPEN,
            carryin => n20824,
            carryout => n20825,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3792__i7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53259\,
            in2 => \_gnd_net_\,
            in3 => \N__53188\,
            lcout => dds0_mclkcnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclkcnt_i7_3792__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16388_2_lut_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53391\,
            in2 => \_gnd_net_\,
            in3 => \N__53217\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclk_297_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__53218\,
            in1 => \N__53364\,
            in2 => \_gnd_net_\,
            in3 => \N__53392\,
            lcout => \DDS_MCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclk_297C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4170_2_lut_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__58193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58030\,
            lcout => OPEN,
            ltout => \n6888_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_72_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__53320\,
            in1 => \N__54175\,
            in2 => \N__53353\,
            in3 => \N__53326\,
            lcout => n21865,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_71_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__63190\,
            in1 => \N__63056\,
            in2 => \N__53338\,
            in3 => \N__57905\,
            lcout => n22027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_75_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__63055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62290\,
            lcout => n22018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_243_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53313\,
            in1 => \N__53301\,
            in2 => \N__53290\,
            in3 => \N__53271\,
            lcout => OPEN,
            ltout => \n12_adj_1685_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_248_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53260\,
            in1 => \N__53244\,
            in2 => \N__53233\,
            in3 => \N__53229\,
            lcout => n21857,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53785\,
            in2 => \_gnd_net_\,
            in3 => \N__53740\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__57078\
        );

    \comm_spi.data_rx_i7_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53781\,
            in1 => \N__53837\,
            in2 => \_gnd_net_\,
            in3 => \N__53739\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i6_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53738\,
            in1 => \N__55132\,
            in2 => \_gnd_net_\,
            in3 => \N__53780\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i5_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53779\,
            in1 => \N__55016\,
            in2 => \_gnd_net_\,
            in3 => \N__53737\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i4_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53736\,
            in1 => \N__62727\,
            in2 => \_gnd_net_\,
            in3 => \N__53778\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i3_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53777\,
            in1 => \N__54878\,
            in2 => \_gnd_net_\,
            in3 => \N__53735\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i2_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53734\,
            in1 => \N__54750\,
            in2 => \_gnd_net_\,
            in3 => \N__53776\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \comm_spi.data_rx_i1_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__53775\,
            in1 => \N__53733\,
            in2 => \_gnd_net_\,
            in3 => \N__54022\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53677\,
            ce => 'H',
            sr => \N__57092\
        );

    \i19760_4_lut_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__63084\,
            in1 => \N__53464\,
            in2 => \N__53455\,
            in3 => \N__61405\,
            lcout => OPEN,
            ltout => \n22321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_1__bdd_4_lut_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__62369\,
            in1 => \N__53446\,
            in2 => \N__53419\,
            in3 => \N__63889\,
            lcout => n23342,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20000_4_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__53409\,
            in1 => \N__58411\,
            in2 => \N__61414\,
            in3 => \N__55558\,
            lcout => n22352,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_299_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54585\,
            in2 => \_gnd_net_\,
            in3 => \N__54444\,
            lcout => n21862,
            ltout => \n21862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i44_4_lut_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__54419\,
            in1 => \N__62368\,
            in2 => \N__54205\,
            in3 => \N__54202\,
            lcout => OPEN,
            ltout => \n22_adj_1725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_294_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__54182\,
            in1 => \N__63083\,
            in2 => \N__54091\,
            in3 => \N__54065\,
            lcout => n12677,
            ltout => \n12677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12759_2_lut_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__63528\,
            in1 => \_gnd_net_\,
            in2 => \N__54088\,
            in3 => \_gnd_net_\,
            lcout => n15482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__63110\,
            in1 => \N__63888\,
            in2 => \_gnd_net_\,
            in3 => \N__63527\,
            lcout => n21895,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i0_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__54037\,
            in1 => \N__62525\,
            in2 => \_gnd_net_\,
            in3 => \N__54021\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i7_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62524\,
            in1 => \N__55884\,
            in2 => \_gnd_net_\,
            in3 => \N__53920\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i6_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53855\,
            in1 => \N__53812\,
            in2 => \_gnd_net_\,
            in3 => \N__62528\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i5_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62523\,
            in1 => \_gnd_net_\,
            in2 => \N__55169\,
            in3 => \N__55105\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i4_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55038\,
            in1 => \N__54991\,
            in2 => \_gnd_net_\,
            in3 => \N__62527\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i3_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__62522\,
            in1 => \_gnd_net_\,
            in2 => \N__62775\,
            in3 => \N__54964\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i2_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__54896\,
            in1 => \N__54850\,
            in2 => \_gnd_net_\,
            in3 => \N__62526\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \comm_buf_4__i1_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__62521\,
            in1 => \N__54769\,
            in2 => \_gnd_net_\,
            in3 => \N__54724\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61942\,
            ce => \N__54694\,
            sr => \N__54688\
        );

    \mux_126_Mux_7_i26_3_lut_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__54676\,
            in1 => \N__59425\,
            in2 => \_gnd_net_\,
            in3 => \N__54657\,
            lcout => OPEN,
            ltout => \n26_adj_1716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19336_4_lut_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__59426\,
            in1 => \N__54628\,
            in2 => \N__54619\,
            in3 => \N__60522\,
            lcout => OPEN,
            ltout => \n22263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_20488_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__59904\,
            in1 => \N__55456\,
            in2 => \N__54616\,
            in3 => \N__60955\,
            lcout => OPEN,
            ltout => \n23420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23420_bdd_4_lut_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__60956\,
            in1 => \N__55999\,
            in2 => \N__55981\,
            in3 => \N__55978\,
            lcout => OPEN,
            ltout => \n23423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_126_Mux_7_i127_3_lut_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55966\,
            in2 => \N__55948\,
            in3 => \N__61409\,
            lcout => OPEN,
            ltout => \comm_buf_1_7_N_559_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__62529\,
            in1 => \N__55899\,
            in2 => \N__55852\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61958\,
            ce => \N__55770\,
            sr => \N__55710\
        );

    \i19746_3_lut_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__55630\,
            in1 => \N__56185\,
            in2 => \_gnd_net_\,
            in3 => \N__58522\,
            lcout => n22356,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23348_bdd_4_lut_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__60516\,
            in1 => \N__55223\,
            in2 => \N__55548\,
            in3 => \N__55510\,
            lcout => n23351,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19335_3_lut_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__60517\,
            in1 => \N__55501\,
            in2 => \_gnd_net_\,
            in3 => \N__55477\,
            lcout => n22262,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20112_2_lut_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__55450\,
            in1 => \_gnd_net_\,
            in2 => \N__59517\,
            in3 => \_gnd_net_\,
            lcout => n22391,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i13_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000101110"
        )
    port map (
            in0 => \N__55227\,
            in1 => \N__55380\,
            in2 => \N__63737\,
            in3 => \N__55288\,
            lcout => buf_dds1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__63643\,
            in1 => \N__56389\,
            in2 => \N__56380\,
            in3 => \N__57730\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61987\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16198_3_lut_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__56532\,
            in1 => \N__56495\,
            in2 => \_gnd_net_\,
            in3 => \N__56478\,
            lcout => n8_adj_1623,
            ltout => \n8_adj_1623_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_358_Mux_5_i15_4_lut_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__63642\,
            in1 => \N__57728\,
            in2 => \N__56383\,
            in3 => \N__56376\,
            lcout => \data_index_9_N_236_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds1_308_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__57729\,
            in1 => \N__63644\,
            in2 => \N__56205\,
            in3 => \N__56257\,
            lcout => trig_dds1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61987\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_298_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__60953\,
            in1 => \N__59900\,
            in2 => \_gnd_net_\,
            in3 => \N__58641\,
            lcout => n21920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19888_4_lut_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000000"
        )
    port map (
            in0 => \N__58642\,
            in1 => \N__60954\,
            in2 => \N__60014\,
            in3 => \N__59400\,
            lcout => OPEN,
            ltout => \n22399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i59_4_lut_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__59401\,
            in1 => \N__56184\,
            in2 => \N__56173\,
            in3 => \N__61401\,
            lcout => n40_adj_1689,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i26_3_lut_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__59497\,
            in1 => \N__56158\,
            in2 => \_gnd_net_\,
            in3 => \N__56133\,
            lcout => n26_adj_1792,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16465_2_lut_3_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__56074\,
            in1 => \N__62646\,
            in2 => \_gnd_net_\,
            in3 => \N__64049\,
            lcout => n14_adj_1611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16456_2_lut_3_lut_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__62056\,
            in1 => \N__62645\,
            in2 => \_gnd_net_\,
            in3 => \N__64048\,
            lcout => n14_adj_1654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i20146_2_lut_4_lut_LC_20_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__64219\,
            in1 => \N__64179\,
            in2 => \N__64168\,
            in3 => \N__64237\,
            lcout => \ADC_VDC.genclk.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i1_LC_20_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64167\,
            in2 => \_gnd_net_\,
            in3 => \N__64220\,
            lcout => \ADC_VDC.genclk.div_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i1C_net\,
            ce => \N__56776\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i20156_2_lut_LC_20_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64162\,
            in2 => \_gnd_net_\,
            in3 => \N__64216\,
            lcout => \ADC_VDC.genclk.n15418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i20142_2_lut_LC_20_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__64217\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__64163\,
            lcout => \ADC_VDC.genclk.n12361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19910_4_lut_LC_20_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__56763\,
            in1 => \N__56751\,
            in2 => \N__56739\,
            in3 => \N__56721\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n22308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i20049_4_lut_LC_20_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57268\,
            in1 => \N__57205\,
            in2 => \N__56710\,
            in3 => \N__56650\,
            lcout => \ADC_VDC.genclk.n22302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_adj_5_LC_20_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56707\,
            in1 => \N__56688\,
            in2 => \N__56677\,
            in3 => \N__56661\,
            lcout => \ADC_VDC.genclk.n27_adj_1483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_adj_3_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56643\,
            in1 => \N__56628\,
            in2 => \N__56617\,
            in3 => \N__56598\,
            lcout => \ADC_VDC.genclk.n28_adj_1481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_adj_4_LC_20_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57261\,
            in1 => \N__57243\,
            in2 => \N__57232\,
            in3 => \N__57216\,
            lcout => \ADC_VDC.genclk.n26_adj_1482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64218\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.genclk.div_state_1__N_1480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_clear_304_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__62450\,
            in1 => \N__63602\,
            in2 => \_gnd_net_\,
            in3 => \N__63072\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61880\,
            ce => \N__56896\,
            sr => \_gnd_net_\
        );

    \i7121_2_lut_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62240\,
            in2 => \_gnd_net_\,
            in3 => \N__63966\,
            lcout => n9837,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20104_2_lut_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56926\,
            in2 => \_gnd_net_\,
            in3 => \N__59420\,
            lcout => n22170,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_144_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__63028\,
            in1 => \N__62242\,
            in2 => \_gnd_net_\,
            in3 => \N__63488\,
            lcout => n12035,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_3_lut_4_lut_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001000100"
        )
    port map (
            in0 => \N__62241\,
            in1 => \N__63027\,
            in2 => \N__58132\,
            in3 => \N__58031\,
            lcout => n7_adj_1687,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_346_Mux_1_i8_3_lut_4_lut_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100000011"
        )
    port map (
            in0 => \N__57907\,
            in1 => \N__56875\,
            in2 => \N__63085\,
            in3 => \N__62296\,
            lcout => n8_adj_1659,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i228_2_lut_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58186\,
            in2 => \_gnd_net_\,
            in3 => \N__58022\,
            lcout => n1373,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_346_Mux_1_i2_3_lut_4_lut_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__62297\,
            in1 => \N__63070\,
            in2 => \N__58205\,
            in3 => \N__57906\,
            lcout => OPEN,
            ltout => \n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23342_bdd_4_lut_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__63071\,
            in1 => \N__63910\,
            in2 => \N__57892\,
            in3 => \N__57889\,
            lcout => OPEN,
            ltout => \n23345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i1_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__57468\,
            in1 => \N__63540\,
            in2 => \N__57367\,
            in3 => \N__57364\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61908\,
            ce => \N__57325\,
            sr => \_gnd_net_\
        );

    \i20047_4_lut_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__62293\,
            in1 => \N__58185\,
            in2 => \N__64029\,
            in3 => \N__57358\,
            lcout => OPEN,
            ltout => \n22340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20168_4_lut_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__57337\,
            in1 => \N__63539\,
            in2 => \N__57328\,
            in3 => \N__63066\,
            lcout => n14_adj_1593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19903_2_lut_3_lut_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110010"
        )
    port map (
            in0 => \N__58035\,
            in1 => \N__63059\,
            in2 => \N__63987\,
            in3 => \_gnd_net_\,
            lcout => n22492,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7001_3_lut_4_lut_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111100100"
        )
    port map (
            in0 => \N__63060\,
            in1 => \N__63908\,
            in2 => \N__57310\,
            in3 => \N__58032\,
            lcout => OPEN,
            ltout => \n9725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_346_Mux_2_i6_4_lut_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__62292\,
            in1 => \N__58187\,
            in2 => \N__57283\,
            in3 => \N__57280\,
            lcout => OPEN,
            ltout => \n6_adj_1657_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__58216\,
            in1 => \N__58237\,
            in2 => \N__58231\,
            in3 => \N__63909\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61921\,
            ce => \N__58225\,
            sr => \N__63617\
        );

    \i1_4_lut_adj_283_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100101100"
        )
    port map (
            in0 => \N__58034\,
            in1 => \N__58192\,
            in2 => \N__63986\,
            in3 => \N__62294\,
            lcout => OPEN,
            ltout => \n26_adj_1597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20171_2_lut_3_lut_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__63058\,
            in1 => \_gnd_net_\,
            in2 => \N__58228\,
            in3 => \N__63541\,
            lcout => n18_adj_1595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_147_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58188\,
            in2 => \_gnd_net_\,
            in3 => \N__62295\,
            lcout => n21908,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_281_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110011"
        )
    port map (
            in0 => \N__63057\,
            in1 => \N__62291\,
            in2 => \N__58206\,
            in3 => \N__58033\,
            lcout => n4_adj_1718,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20087_2_lut_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58915\,
            in2 => \_gnd_net_\,
            in3 => \N__57958\,
            lcout => n22642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_5_i127_3_lut_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57937\,
            in1 => \N__58318\,
            in2 => \_gnd_net_\,
            in3 => \N__61406\,
            lcout => \comm_buf_0_7_N_543_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_300_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011111011"
        )
    port map (
            in0 => \N__59421\,
            in1 => \N__61034\,
            in2 => \N__60044\,
            in3 => \N__60499\,
            lcout => n48,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19784_2_lut_3_lut_4_lut_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__58653\,
            in1 => \N__58492\,
            in2 => \N__60043\,
            in3 => \N__61033\,
            lcout => n22365,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19803_3_lut_4_lut_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__61035\,
            in1 => \N__58654\,
            in2 => \N__58511\,
            in3 => \N__59423\,
            lcout => OPEN,
            ltout => \n22364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20094_4_lut_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__58429\,
            in1 => \N__61374\,
            in2 => \N__58423\,
            in3 => \N__60501\,
            lcout => OPEN,
            ltout => \n22370_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19802_4_lut_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__61375\,
            in1 => \N__58420\,
            in2 => \N__58414\,
            in3 => \N__58407\,
            lcout => n22368,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_185_i9_2_lut_3_lut_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__59422\,
            in1 => \N__59954\,
            in2 => \_gnd_net_\,
            in3 => \N__60500\,
            lcout => n9_adj_1507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23492_bdd_4_lut_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__61036\,
            in1 => \N__58348\,
            in2 => \N__58330\,
            in3 => \N__60721\,
            lcout => n23495,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19755_2_lut_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58312\,
            in2 => \_gnd_net_\,
            in3 => \N__59424\,
            lcout => n22316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n23456_bdd_4_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__60093\,
            in1 => \N__58300\,
            in2 => \N__58291\,
            in3 => \N__59566\,
            lcout => OPEN,
            ltout => \n23459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1661462_i1_3_lut_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58276\,
            in2 => \N__58258\,
            in3 => \N__61020\,
            lcout => OPEN,
            ltout => \n30_adj_1793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_3_i127_3_lut_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58255\,
            in2 => \N__61417\,
            in3 => \N__61410\,
            lcout => \comm_buf_0_7_N_543_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_5_i28_4_lut_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001001000000"
        )
    port map (
            in0 => \N__60601\,
            in1 => \N__59406\,
            in2 => \N__61102\,
            in3 => \N__61075\,
            lcout => OPEN,
            ltout => \n28_adj_1775_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__60676\,
            in1 => \N__60092\,
            in2 => \N__61060\,
            in3 => \N__61019\,
            lcout => n23492,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_125_Mux_5_i25_4_lut_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__60600\,
            in1 => \N__59405\,
            in2 => \N__60712\,
            in3 => \N__60697\,
            lcout => n25_adj_1774,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_20508_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__60602\,
            in1 => \N__60064\,
            in2 => \N__59584\,
            in3 => \N__59572\,
            lcout => n23456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19937_2_lut_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59560\,
            in2 => \_gnd_net_\,
            in3 => \N__59501\,
            lcout => n22313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19751_2_lut_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59542\,
            in2 => \_gnd_net_\,
            in3 => \N__59407\,
            lcout => n22300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20099_2_lut_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59527\,
            in2 => \_gnd_net_\,
            in3 => \N__59496\,
            lcout => n22649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_LC_22_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__64902\,
            in1 => \N__64341\,
            in2 => \N__64984\,
            in3 => \N__64302\,
            lcout => \ADC_VDC.genclk.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_LC_22_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__64917\,
            in1 => \N__64359\,
            in2 => \N__64270\,
            in3 => \N__64947\,
            lcout => \ADC_VDC.genclk.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i20011_4_lut_LC_22_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__64284\,
            in1 => \N__64377\,
            in2 => \N__64327\,
            in3 => \N__64392\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n22305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19909_4_lut_LC_22_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__64138\,
            in1 => \N__64252\,
            in2 => \N__64246\,
            in3 => \N__64243\,
            lcout => \ADC_VDC.genclk.n22303\,
            ltout => \ADC_VDC.genclk.n22303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i0_LC_22_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__64161\,
            in1 => \N__64228\,
            in2 => \N__64189\,
            in3 => \N__64186\,
            lcout => \ADC_VDC.genclk.div_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_LC_22_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__64887\,
            in1 => \N__64962\,
            in2 => \N__64498\,
            in3 => \N__64932\,
            lcout => \ADC_VDC.genclk.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_response_305_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000110100"
        )
    port map (
            in0 => \N__64025\,
            in1 => \N__63491\,
            in2 => \N__62633\,
            in3 => \N__63077\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61924\,
            ce => \N__62803\,
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010000"
        )
    port map (
            in0 => \N__63959\,
            in1 => \N__63722\,
            in2 => \N__63205\,
            in3 => \N__63074\,
            lcout => n12045,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i3_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__62780\,
            in1 => \N__62602\,
            in2 => \_gnd_net_\,
            in3 => \N__62113\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__61976\,
            ce => \N__61437\,
            sr => \N__64416\
        );

    \ADC_VDC.genclk.t0off_i0_LC_23_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64393\,
            in2 => \_gnd_net_\,
            in3 => \N__64381\,
            lcout => \ADC_VDC.genclk.t0off_0\,
            ltout => OPEN,
            carryin => \bfn_23_5_0_\,
            carryout => \ADC_VDC.genclk.n20736\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i1_LC_23_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64378\,
            in2 => \N__64848\,
            in3 => \N__64366\,
            lcout => \ADC_VDC.genclk.t0off_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20736\,
            carryout => \ADC_VDC.genclk.n20737\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i2_LC_23_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64795\,
            in2 => \N__64363\,
            in3 => \N__64345\,
            lcout => \ADC_VDC.genclk.t0off_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20737\,
            carryout => \ADC_VDC.genclk.n20738\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i3_LC_23_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64342\,
            in2 => \N__64849\,
            in3 => \N__64330\,
            lcout => \ADC_VDC.genclk.t0off_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20738\,
            carryout => \ADC_VDC.genclk.n20739\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i4_LC_23_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64799\,
            in2 => \N__64326\,
            in3 => \N__64306\,
            lcout => \ADC_VDC.genclk.t0off_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20739\,
            carryout => \ADC_VDC.genclk.n20740\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i5_LC_23_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64303\,
            in2 => \N__64850\,
            in3 => \N__64291\,
            lcout => \ADC_VDC.genclk.t0off_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20740\,
            carryout => \ADC_VDC.genclk.n20741\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i6_LC_23_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64803\,
            in2 => \N__64288\,
            in3 => \N__64273\,
            lcout => \ADC_VDC.genclk.t0off_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20741\,
            carryout => \ADC_VDC.genclk.n20742\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i7_LC_23_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64269\,
            in2 => \N__64851\,
            in3 => \N__64255\,
            lcout => \ADC_VDC.genclk.t0off_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20742\,
            carryout => \ADC_VDC.genclk.n20743\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__64479\,
            sr => \N__64459\
        );

    \ADC_VDC.genclk.t0off_i8_LC_23_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64980\,
            in2 => \N__64730\,
            in3 => \N__64966\,
            lcout => \ADC_VDC.genclk.t0off_8\,
            ltout => OPEN,
            carryin => \bfn_23_6_0_\,
            carryout => \ADC_VDC.genclk.n20744\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i9_LC_23_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64963\,
            in2 => \N__64733\,
            in3 => \N__64951\,
            lcout => \ADC_VDC.genclk.t0off_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20744\,
            carryout => \ADC_VDC.genclk.n20745\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i10_LC_23_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64948\,
            in2 => \N__64727\,
            in3 => \N__64936\,
            lcout => \ADC_VDC.genclk.t0off_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20745\,
            carryout => \ADC_VDC.genclk.n20746\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i11_LC_23_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64933\,
            in2 => \N__64731\,
            in3 => \N__64921\,
            lcout => \ADC_VDC.genclk.t0off_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20746\,
            carryout => \ADC_VDC.genclk.n20747\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i12_LC_23_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64918\,
            in2 => \N__64728\,
            in3 => \N__64906\,
            lcout => \ADC_VDC.genclk.t0off_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20747\,
            carryout => \ADC_VDC.genclk.n20748\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i13_LC_23_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64903\,
            in2 => \N__64732\,
            in3 => \N__64891\,
            lcout => \ADC_VDC.genclk.t0off_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20748\,
            carryout => \ADC_VDC.genclk.n20749\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i14_LC_23_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64888\,
            in2 => \N__64729\,
            in3 => \N__64876\,
            lcout => \ADC_VDC.genclk.t0off_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n20749\,
            carryout => \ADC_VDC.genclk.n20750\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );

    \ADC_VDC.genclk.t0off_i15_LC_23_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__64666\,
            in1 => \N__64497\,
            in2 => \_gnd_net_\,
            in3 => \N__64501\,
            lcout => \ADC_VDC.genclk.t0off_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__64483\,
            sr => \N__64458\
        );
end \INTERFACE\;
