-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 28 2024 17:12:44

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zim" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zim
entity zim is
port (
    VAC_DRDY : in std_logic;
    IAC_FLT1 : out std_logic;
    DDS_SCK : out std_logic;
    ICE_IOR_166 : in std_logic;
    ICE_IOR_119 : in std_logic;
    DDS_MOSI : out std_logic;
    VAC_MISO : in std_logic;
    DDS_MOSI1 : out std_logic;
    ICE_IOR_146 : in std_logic;
    VDC_CLK : out std_logic;
    ICE_IOT_222 : in std_logic;
    IAC_CS : out std_logic;
    ICE_IOL_18B : in std_logic;
    ICE_IOL_13A : in std_logic;
    ICE_IOB_81 : in std_logic;
    VAC_OSR1 : out std_logic;
    IAC_MOSI : out std_logic;
    DDS_CS1 : out std_logic;
    ICE_IOL_4B : in std_logic;
    ICE_IOB_94 : in std_logic;
    VAC_CS : out std_logic;
    VAC_CLK : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    ICE_IOR_167 : in std_logic;
    ICE_IOR_118 : in std_logic;
    RTD_SDO : in std_logic;
    IAC_OSR0 : out std_logic;
    VDC_SCLK : out std_logic;
    VAC_FLT1 : out std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_IOR_165 : in std_logic;
    ICE_IOR_147 : in std_logic;
    ICE_IOL_14A : in std_logic;
    ICE_IOL_13B : in std_logic;
    ICE_IOB_91 : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_RNG_0 : out std_logic;
    VDC_RNG0 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    ICE_IOR_152 : in std_logic;
    ICE_IOL_12A : in std_logic;
    RTD_DRDY : in std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_IOT_177 : in std_logic;
    ICE_IOR_141 : in std_logic;
    ICE_IOB_102 : in std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    IAC_MISO : in std_logic;
    VAC_OSR0 : out std_logic;
    VAC_MOSI : out std_logic;
    TEST_LED : out std_logic;
    ICE_IOR_148 : in std_logic;
    STAT_COMM : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_IOR_161 : in std_logic;
    ICE_IOB_95 : in std_logic;
    ICE_IOB_82 : in std_logic;
    ICE_IOB_104 : in std_logic;
    IAC_CLK : out std_logic;
    DDS_CS : out std_logic;
    SELIRNG0 : out std_logic;
    RTD_SDI : out std_logic;
    ICE_IOT_221 : in std_logic;
    ICE_IOT_197 : in std_logic;
    DDS_MCLK : out std_logic;
    RTD_SCLK : out std_logic;
    RTD_CS : out std_logic;
    ICE_IOR_137 : in std_logic;
    IAC_OSR1 : out std_logic;
    VAC_FLT0 : out std_logic;
    ICE_IOR_144 : in std_logic;
    ICE_IOR_128 : in std_logic;
    ICE_GPMO_1 : in std_logic;
    IAC_SCLK : out std_logic;
    EIS_SYNCCLK : in std_logic;
    ICE_IOR_139 : in std_logic;
    ICE_IOL_4A : in std_logic;
    VAC_SCLK : out std_logic;
    THERMOSTAT : in std_logic;
    ICE_IOR_164 : in std_logic;
    ICE_IOB_103 : in std_logic;
    OUT_SYNCCLK : out std_logic;
    AMPV_POW : out std_logic;
    VDC_SDO : in std_logic;
    ICE_IOT_174 : in std_logic;
    ICE_IOR_140 : in std_logic;
    ICE_IOB_96 : in std_logic;
    CONT_SD : out std_logic;
    AC_ADC_SYNC : out std_logic;
    SELIRNG1 : out std_logic;
    ICE_IOL_12B : in std_logic;
    ICE_IOR_160 : in std_logic;
    ICE_IOR_136 : in std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_IOT_198 : in std_logic;
    ICE_IOT_173 : in std_logic;
    IAC_DRDY : in std_logic;
    ICE_IOT_178 : in std_logic;
    ICE_IOR_138 : in std_logic;
    ICE_IOR_120 : in std_logic;
    IAC_FLT0 : out std_logic;
    DDS_SCK1 : out std_logic);
end zim;

-- Architecture of zim
-- View name is \INTERFACE\
architecture \INTERFACE\ of zim is

signal \N__59184\ : std_logic;
signal \N__59183\ : std_logic;
signal \N__59182\ : std_logic;
signal \N__59175\ : std_logic;
signal \N__59174\ : std_logic;
signal \N__59173\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59164\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59156\ : std_logic;
signal \N__59155\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59146\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59137\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59129\ : std_logic;
signal \N__59128\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59110\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59094\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59092\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59084\ : std_logic;
signal \N__59083\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__59067\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59065\ : std_logic;
signal \N__59058\ : std_logic;
signal \N__59057\ : std_logic;
signal \N__59056\ : std_logic;
signal \N__59049\ : std_logic;
signal \N__59048\ : std_logic;
signal \N__59047\ : std_logic;
signal \N__59040\ : std_logic;
signal \N__59039\ : std_logic;
signal \N__59038\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59030\ : std_logic;
signal \N__59029\ : std_logic;
signal \N__59022\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59020\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59012\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59004\ : std_logic;
signal \N__59003\ : std_logic;
signal \N__59002\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58994\ : std_logic;
signal \N__58993\ : std_logic;
signal \N__58986\ : std_logic;
signal \N__58985\ : std_logic;
signal \N__58984\ : std_logic;
signal \N__58977\ : std_logic;
signal \N__58976\ : std_logic;
signal \N__58975\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58967\ : std_logic;
signal \N__58966\ : std_logic;
signal \N__58959\ : std_logic;
signal \N__58958\ : std_logic;
signal \N__58957\ : std_logic;
signal \N__58950\ : std_logic;
signal \N__58949\ : std_logic;
signal \N__58948\ : std_logic;
signal \N__58941\ : std_logic;
signal \N__58940\ : std_logic;
signal \N__58939\ : std_logic;
signal \N__58932\ : std_logic;
signal \N__58931\ : std_logic;
signal \N__58930\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58922\ : std_logic;
signal \N__58921\ : std_logic;
signal \N__58914\ : std_logic;
signal \N__58913\ : std_logic;
signal \N__58912\ : std_logic;
signal \N__58905\ : std_logic;
signal \N__58904\ : std_logic;
signal \N__58903\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58895\ : std_logic;
signal \N__58894\ : std_logic;
signal \N__58887\ : std_logic;
signal \N__58886\ : std_logic;
signal \N__58885\ : std_logic;
signal \N__58878\ : std_logic;
signal \N__58877\ : std_logic;
signal \N__58876\ : std_logic;
signal \N__58869\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58867\ : std_logic;
signal \N__58860\ : std_logic;
signal \N__58859\ : std_logic;
signal \N__58858\ : std_logic;
signal \N__58851\ : std_logic;
signal \N__58850\ : std_logic;
signal \N__58849\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58841\ : std_logic;
signal \N__58840\ : std_logic;
signal \N__58833\ : std_logic;
signal \N__58832\ : std_logic;
signal \N__58831\ : std_logic;
signal \N__58824\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58822\ : std_logic;
signal \N__58815\ : std_logic;
signal \N__58814\ : std_logic;
signal \N__58813\ : std_logic;
signal \N__58806\ : std_logic;
signal \N__58805\ : std_logic;
signal \N__58804\ : std_logic;
signal \N__58797\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58795\ : std_logic;
signal \N__58788\ : std_logic;
signal \N__58787\ : std_logic;
signal \N__58786\ : std_logic;
signal \N__58779\ : std_logic;
signal \N__58778\ : std_logic;
signal \N__58777\ : std_logic;
signal \N__58770\ : std_logic;
signal \N__58769\ : std_logic;
signal \N__58768\ : std_logic;
signal \N__58761\ : std_logic;
signal \N__58760\ : std_logic;
signal \N__58759\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58751\ : std_logic;
signal \N__58750\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58742\ : std_logic;
signal \N__58741\ : std_logic;
signal \N__58734\ : std_logic;
signal \N__58733\ : std_logic;
signal \N__58732\ : std_logic;
signal \N__58725\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58723\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58715\ : std_logic;
signal \N__58714\ : std_logic;
signal \N__58707\ : std_logic;
signal \N__58706\ : std_logic;
signal \N__58705\ : std_logic;
signal \N__58698\ : std_logic;
signal \N__58697\ : std_logic;
signal \N__58696\ : std_logic;
signal \N__58689\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58687\ : std_logic;
signal \N__58680\ : std_logic;
signal \N__58679\ : std_logic;
signal \N__58678\ : std_logic;
signal \N__58671\ : std_logic;
signal \N__58670\ : std_logic;
signal \N__58669\ : std_logic;
signal \N__58662\ : std_logic;
signal \N__58661\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58653\ : std_logic;
signal \N__58652\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58644\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58642\ : std_logic;
signal \N__58635\ : std_logic;
signal \N__58634\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58625\ : std_logic;
signal \N__58624\ : std_logic;
signal \N__58617\ : std_logic;
signal \N__58616\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58608\ : std_logic;
signal \N__58607\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58598\ : std_logic;
signal \N__58597\ : std_logic;
signal \N__58590\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58588\ : std_logic;
signal \N__58581\ : std_logic;
signal \N__58580\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58572\ : std_logic;
signal \N__58571\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58563\ : std_logic;
signal \N__58562\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58554\ : std_logic;
signal \N__58553\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58545\ : std_logic;
signal \N__58544\ : std_logic;
signal \N__58543\ : std_logic;
signal \N__58536\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58527\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58518\ : std_logic;
signal \N__58517\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58509\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58489\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58481\ : std_logic;
signal \N__58480\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58472\ : std_logic;
signal \N__58471\ : std_logic;
signal \N__58464\ : std_logic;
signal \N__58463\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58454\ : std_logic;
signal \N__58453\ : std_logic;
signal \N__58446\ : std_logic;
signal \N__58445\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58437\ : std_logic;
signal \N__58436\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58427\ : std_logic;
signal \N__58426\ : std_logic;
signal \N__58419\ : std_logic;
signal \N__58418\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58410\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58401\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58391\ : std_logic;
signal \N__58390\ : std_logic;
signal \N__58383\ : std_logic;
signal \N__58382\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58374\ : std_logic;
signal \N__58373\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58364\ : std_logic;
signal \N__58363\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58355\ : std_logic;
signal \N__58354\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58346\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58338\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58329\ : std_logic;
signal \N__58328\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58320\ : std_logic;
signal \N__58319\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58311\ : std_logic;
signal \N__58310\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58302\ : std_logic;
signal \N__58301\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58293\ : std_logic;
signal \N__58292\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58283\ : std_logic;
signal \N__58282\ : std_logic;
signal \N__58275\ : std_logic;
signal \N__58274\ : std_logic;
signal \N__58273\ : std_logic;
signal \N__58266\ : std_logic;
signal \N__58265\ : std_logic;
signal \N__58264\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58244\ : std_logic;
signal \N__58241\ : std_logic;
signal \N__58238\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58234\ : std_logic;
signal \N__58231\ : std_logic;
signal \N__58228\ : std_logic;
signal \N__58225\ : std_logic;
signal \N__58224\ : std_logic;
signal \N__58221\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58215\ : std_logic;
signal \N__58208\ : std_logic;
signal \N__58207\ : std_logic;
signal \N__58204\ : std_logic;
signal \N__58201\ : std_logic;
signal \N__58198\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58192\ : std_logic;
signal \N__58189\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58178\ : std_logic;
signal \N__58177\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58171\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58163\ : std_logic;
signal \N__58160\ : std_logic;
signal \N__58157\ : std_logic;
signal \N__58154\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58152\ : std_logic;
signal \N__58149\ : std_logic;
signal \N__58146\ : std_logic;
signal \N__58143\ : std_logic;
signal \N__58136\ : std_logic;
signal \N__58135\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58128\ : std_logic;
signal \N__58125\ : std_logic;
signal \N__58122\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58116\ : std_logic;
signal \N__58113\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58103\ : std_logic;
signal \N__58100\ : std_logic;
signal \N__58097\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58091\ : std_logic;
signal \N__58088\ : std_logic;
signal \N__58085\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58078\ : std_logic;
signal \N__58073\ : std_logic;
signal \N__58070\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58064\ : std_logic;
signal \N__58061\ : std_logic;
signal \N__58058\ : std_logic;
signal \N__58055\ : std_logic;
signal \N__58054\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58048\ : std_logic;
signal \N__58045\ : std_logic;
signal \N__58042\ : std_logic;
signal \N__58041\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58035\ : std_logic;
signal \N__58032\ : std_logic;
signal \N__58031\ : std_logic;
signal \N__58030\ : std_logic;
signal \N__58025\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58019\ : std_logic;
signal \N__58016\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58006\ : std_logic;
signal \N__58001\ : std_logic;
signal \N__57998\ : std_logic;
signal \N__57995\ : std_logic;
signal \N__57992\ : std_logic;
signal \N__57989\ : std_logic;
signal \N__57986\ : std_logic;
signal \N__57983\ : std_logic;
signal \N__57982\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57980\ : std_logic;
signal \N__57979\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57977\ : std_logic;
signal \N__57976\ : std_logic;
signal \N__57975\ : std_logic;
signal \N__57974\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57972\ : std_logic;
signal \N__57971\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57968\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57965\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57962\ : std_logic;
signal \N__57961\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57956\ : std_logic;
signal \N__57955\ : std_logic;
signal \N__57954\ : std_logic;
signal \N__57953\ : std_logic;
signal \N__57952\ : std_logic;
signal \N__57951\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57948\ : std_logic;
signal \N__57947\ : std_logic;
signal \N__57946\ : std_logic;
signal \N__57945\ : std_logic;
signal \N__57944\ : std_logic;
signal \N__57943\ : std_logic;
signal \N__57942\ : std_logic;
signal \N__57941\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57939\ : std_logic;
signal \N__57938\ : std_logic;
signal \N__57937\ : std_logic;
signal \N__57936\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57934\ : std_logic;
signal \N__57933\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57930\ : std_logic;
signal \N__57929\ : std_logic;
signal \N__57928\ : std_logic;
signal \N__57927\ : std_logic;
signal \N__57926\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57924\ : std_logic;
signal \N__57923\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57921\ : std_logic;
signal \N__57920\ : std_logic;
signal \N__57919\ : std_logic;
signal \N__57918\ : std_logic;
signal \N__57917\ : std_logic;
signal \N__57916\ : std_logic;
signal \N__57915\ : std_logic;
signal \N__57914\ : std_logic;
signal \N__57913\ : std_logic;
signal \N__57912\ : std_logic;
signal \N__57911\ : std_logic;
signal \N__57910\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57908\ : std_logic;
signal \N__57907\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57904\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57902\ : std_logic;
signal \N__57901\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57899\ : std_logic;
signal \N__57898\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57895\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57893\ : std_logic;
signal \N__57892\ : std_logic;
signal \N__57891\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57888\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57885\ : std_logic;
signal \N__57884\ : std_logic;
signal \N__57883\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57881\ : std_logic;
signal \N__57880\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57875\ : std_logic;
signal \N__57874\ : std_logic;
signal \N__57873\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57870\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57868\ : std_logic;
signal \N__57867\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57865\ : std_logic;
signal \N__57864\ : std_logic;
signal \N__57863\ : std_logic;
signal \N__57862\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57857\ : std_logic;
signal \N__57856\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57854\ : std_logic;
signal \N__57853\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57851\ : std_logic;
signal \N__57850\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57848\ : std_logic;
signal \N__57847\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57845\ : std_logic;
signal \N__57844\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57842\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57839\ : std_logic;
signal \N__57838\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57836\ : std_logic;
signal \N__57835\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57832\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57829\ : std_logic;
signal \N__57828\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57826\ : std_logic;
signal \N__57825\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57822\ : std_logic;
signal \N__57821\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57818\ : std_logic;
signal \N__57817\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57815\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57812\ : std_logic;
signal \N__57811\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57809\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57807\ : std_logic;
signal \N__57806\ : std_logic;
signal \N__57805\ : std_logic;
signal \N__57804\ : std_logic;
signal \N__57443\ : std_logic;
signal \N__57440\ : std_logic;
signal \N__57437\ : std_logic;
signal \N__57434\ : std_logic;
signal \N__57431\ : std_logic;
signal \N__57428\ : std_logic;
signal \N__57425\ : std_logic;
signal \N__57424\ : std_logic;
signal \N__57423\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57418\ : std_logic;
signal \N__57415\ : std_logic;
signal \N__57414\ : std_logic;
signal \N__57411\ : std_logic;
signal \N__57410\ : std_logic;
signal \N__57395\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57391\ : std_logic;
signal \N__57390\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57385\ : std_logic;
signal \N__57384\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57382\ : std_logic;
signal \N__57381\ : std_logic;
signal \N__57380\ : std_logic;
signal \N__57379\ : std_logic;
signal \N__57376\ : std_logic;
signal \N__57375\ : std_logic;
signal \N__57374\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57369\ : std_logic;
signal \N__57366\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57358\ : std_logic;
signal \N__57357\ : std_logic;
signal \N__57354\ : std_logic;
signal \N__57353\ : std_logic;
signal \N__57350\ : std_logic;
signal \N__57347\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57342\ : std_logic;
signal \N__57339\ : std_logic;
signal \N__57338\ : std_logic;
signal \N__57335\ : std_logic;
signal \N__57334\ : std_logic;
signal \N__57331\ : std_logic;
signal \N__57328\ : std_logic;
signal \N__57327\ : std_logic;
signal \N__57326\ : std_logic;
signal \N__57325\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57321\ : std_logic;
signal \N__57320\ : std_logic;
signal \N__57319\ : std_logic;
signal \N__57318\ : std_logic;
signal \N__57301\ : std_logic;
signal \N__57286\ : std_logic;
signal \N__57283\ : std_logic;
signal \N__57266\ : std_logic;
signal \N__57263\ : std_logic;
signal \N__57260\ : std_logic;
signal \N__57259\ : std_logic;
signal \N__57256\ : std_logic;
signal \N__57255\ : std_logic;
signal \N__57252\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57248\ : std_logic;
signal \N__57245\ : std_logic;
signal \N__57242\ : std_logic;
signal \N__57239\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57237\ : std_logic;
signal \N__57236\ : std_logic;
signal \N__57233\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57227\ : std_logic;
signal \N__57222\ : std_logic;
signal \N__57219\ : std_logic;
signal \N__57204\ : std_logic;
signal \N__57197\ : std_logic;
signal \N__57194\ : std_logic;
signal \N__57191\ : std_logic;
signal \N__57188\ : std_logic;
signal \N__57187\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57185\ : std_logic;
signal \N__57182\ : std_logic;
signal \N__57179\ : std_logic;
signal \N__57174\ : std_logic;
signal \N__57171\ : std_logic;
signal \N__57168\ : std_logic;
signal \N__57167\ : std_logic;
signal \N__57158\ : std_logic;
signal \N__57155\ : std_logic;
signal \N__57152\ : std_logic;
signal \N__57149\ : std_logic;
signal \N__57148\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57144\ : std_logic;
signal \N__57141\ : std_logic;
signal \N__57138\ : std_logic;
signal \N__57133\ : std_logic;
signal \N__57130\ : std_logic;
signal \N__57121\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57112\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57106\ : std_logic;
signal \N__57103\ : std_logic;
signal \N__57100\ : std_logic;
signal \N__57093\ : std_logic;
signal \N__57080\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57070\ : std_logic;
signal \N__57067\ : std_logic;
signal \N__57062\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57058\ : std_logic;
signal \N__57055\ : std_logic;
signal \N__57052\ : std_logic;
signal \N__57051\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57049\ : std_logic;
signal \N__57044\ : std_logic;
signal \N__57041\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57037\ : std_logic;
signal \N__57036\ : std_logic;
signal \N__57035\ : std_logic;
signal \N__57032\ : std_logic;
signal \N__57027\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__57017\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57013\ : std_logic;
signal \N__57012\ : std_logic;
signal \N__57009\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__56999\ : std_logic;
signal \N__56998\ : std_logic;
signal \N__56997\ : std_logic;
signal \N__56996\ : std_logic;
signal \N__56995\ : std_logic;
signal \N__56992\ : std_logic;
signal \N__56991\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56987\ : std_logic;
signal \N__56984\ : std_logic;
signal \N__56983\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56975\ : std_logic;
signal \N__56972\ : std_logic;
signal \N__56969\ : std_logic;
signal \N__56966\ : std_logic;
signal \N__56963\ : std_logic;
signal \N__56960\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56954\ : std_logic;
signal \N__56951\ : std_logic;
signal \N__56948\ : std_logic;
signal \N__56945\ : std_logic;
signal \N__56942\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56936\ : std_logic;
signal \N__56931\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56919\ : std_logic;
signal \N__56918\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56912\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56907\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56892\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56883\ : std_logic;
signal \N__56880\ : std_logic;
signal \N__56877\ : std_logic;
signal \N__56858\ : std_logic;
signal \N__56855\ : std_logic;
signal \N__56854\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56852\ : std_logic;
signal \N__56849\ : std_logic;
signal \N__56846\ : std_logic;
signal \N__56845\ : std_logic;
signal \N__56844\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56842\ : std_logic;
signal \N__56841\ : std_logic;
signal \N__56838\ : std_logic;
signal \N__56837\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56818\ : std_logic;
signal \N__56817\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56808\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56795\ : std_logic;
signal \N__56792\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56777\ : std_logic;
signal \N__56776\ : std_logic;
signal \N__56775\ : std_logic;
signal \N__56772\ : std_logic;
signal \N__56767\ : std_logic;
signal \N__56764\ : std_logic;
signal \N__56761\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56755\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56750\ : std_logic;
signal \N__56749\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56747\ : std_logic;
signal \N__56746\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56744\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56737\ : std_logic;
signal \N__56732\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56724\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56716\ : std_logic;
signal \N__56713\ : std_logic;
signal \N__56706\ : std_logic;
signal \N__56703\ : std_logic;
signal \N__56698\ : std_logic;
signal \N__56695\ : std_logic;
signal \N__56684\ : std_logic;
signal \N__56675\ : std_logic;
signal \N__56672\ : std_logic;
signal \N__56667\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56633\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56628\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56622\ : std_logic;
signal \N__56619\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56611\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56605\ : std_logic;
signal \N__56600\ : std_logic;
signal \N__56597\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56591\ : std_logic;
signal \N__56588\ : std_logic;
signal \N__56585\ : std_logic;
signal \N__56584\ : std_logic;
signal \N__56581\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56577\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56549\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56542\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56535\ : std_logic;
signal \N__56530\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56524\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56516\ : std_logic;
signal \N__56513\ : std_logic;
signal \N__56510\ : std_logic;
signal \N__56507\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56505\ : std_logic;
signal \N__56502\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56496\ : std_logic;
signal \N__56489\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56475\ : std_logic;
signal \N__56470\ : std_logic;
signal \N__56467\ : std_logic;
signal \N__56464\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56449\ : std_logic;
signal \N__56444\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56438\ : std_logic;
signal \N__56435\ : std_logic;
signal \N__56432\ : std_logic;
signal \N__56429\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56425\ : std_logic;
signal \N__56422\ : std_logic;
signal \N__56419\ : std_logic;
signal \N__56414\ : std_logic;
signal \N__56411\ : std_logic;
signal \N__56408\ : std_logic;
signal \N__56405\ : std_logic;
signal \N__56402\ : std_logic;
signal \N__56399\ : std_logic;
signal \N__56396\ : std_logic;
signal \N__56395\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56385\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56377\ : std_logic;
signal \N__56374\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56372\ : std_logic;
signal \N__56371\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56369\ : std_logic;
signal \N__56368\ : std_logic;
signal \N__56367\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56340\ : std_logic;
signal \N__56339\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56337\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56332\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56330\ : std_logic;
signal \N__56329\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56320\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56318\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56314\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56310\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56306\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56303\ : std_logic;
signal \N__56302\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56300\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56282\ : std_logic;
signal \N__56281\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56264\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56237\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56231\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56216\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56210\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56187\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56185\ : std_logic;
signal \N__56184\ : std_logic;
signal \N__56183\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56177\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56171\ : std_logic;
signal \N__56168\ : std_logic;
signal \N__56167\ : std_logic;
signal \N__56166\ : std_logic;
signal \N__56163\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56159\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56137\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56123\ : std_logic;
signal \N__56120\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56094\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56072\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56061\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56032\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56009\ : std_logic;
signal \N__56008\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56006\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55988\ : std_logic;
signal \N__55985\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55970\ : std_logic;
signal \N__55967\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55948\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55935\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55929\ : std_logic;
signal \N__55924\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55914\ : std_logic;
signal \N__55909\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55881\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55857\ : std_logic;
signal \N__55850\ : std_logic;
signal \N__55847\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55803\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55788\ : std_logic;
signal \N__55781\ : std_logic;
signal \N__55770\ : std_logic;
signal \N__55755\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55735\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55703\ : std_logic;
signal \N__55700\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55691\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55684\ : std_logic;
signal \N__55681\ : std_logic;
signal \N__55678\ : std_logic;
signal \N__55673\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55658\ : std_logic;
signal \N__55655\ : std_logic;
signal \N__55654\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55636\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55624\ : std_logic;
signal \N__55619\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55607\ : std_logic;
signal \N__55604\ : std_logic;
signal \N__55601\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55583\ : std_logic;
signal \N__55580\ : std_logic;
signal \N__55577\ : std_logic;
signal \N__55574\ : std_logic;
signal \N__55571\ : std_logic;
signal \N__55568\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55562\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55547\ : std_logic;
signal \N__55544\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55520\ : std_logic;
signal \N__55517\ : std_logic;
signal \N__55514\ : std_logic;
signal \N__55511\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55498\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55484\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55457\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55440\ : std_logic;
signal \N__55437\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55411\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55397\ : std_logic;
signal \N__55394\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55390\ : std_logic;
signal \N__55387\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55373\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55367\ : std_logic;
signal \N__55366\ : std_logic;
signal \N__55363\ : std_logic;
signal \N__55360\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55354\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55343\ : std_logic;
signal \N__55340\ : std_logic;
signal \N__55339\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55318\ : std_logic;
signal \N__55315\ : std_logic;
signal \N__55312\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55308\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55267\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55259\ : std_logic;
signal \N__55256\ : std_logic;
signal \N__55253\ : std_logic;
signal \N__55250\ : std_logic;
signal \N__55247\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55226\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55201\ : std_logic;
signal \N__55198\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55153\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55135\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55112\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55106\ : std_logic;
signal \N__55103\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55094\ : std_logic;
signal \N__55091\ : std_logic;
signal \N__55088\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55052\ : std_logic;
signal \N__55049\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55043\ : std_logic;
signal \N__55040\ : std_logic;
signal \N__55039\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55024\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55008\ : std_logic;
signal \N__55003\ : std_logic;
signal \N__55000\ : std_logic;
signal \N__54997\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54989\ : std_logic;
signal \N__54986\ : std_logic;
signal \N__54983\ : std_logic;
signal \N__54982\ : std_logic;
signal \N__54981\ : std_logic;
signal \N__54978\ : std_logic;
signal \N__54977\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54974\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54972\ : std_logic;
signal \N__54971\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54966\ : std_logic;
signal \N__54965\ : std_logic;
signal \N__54964\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54962\ : std_logic;
signal \N__54961\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54954\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54949\ : std_logic;
signal \N__54948\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54945\ : std_logic;
signal \N__54932\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54913\ : std_logic;
signal \N__54912\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54907\ : std_logic;
signal \N__54904\ : std_logic;
signal \N__54903\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54901\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54899\ : std_logic;
signal \N__54896\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54892\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54870\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54867\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54846\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54830\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54824\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54818\ : std_logic;
signal \N__54811\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54809\ : std_logic;
signal \N__54808\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54766\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54763\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54735\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54722\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54717\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54707\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54705\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54661\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54655\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54641\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54637\ : std_logic;
signal \N__54636\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54629\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54621\ : std_logic;
signal \N__54616\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54605\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54560\ : std_logic;
signal \N__54559\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54548\ : std_logic;
signal \N__54545\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54537\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54530\ : std_logic;
signal \N__54529\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54496\ : std_logic;
signal \N__54493\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54479\ : std_logic;
signal \N__54476\ : std_logic;
signal \N__54471\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54463\ : std_logic;
signal \N__54456\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54425\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54382\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54378\ : std_logic;
signal \N__54375\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54372\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54369\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54356\ : std_logic;
signal \N__54353\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54344\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54330\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54319\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54291\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54273\ : std_logic;
signal \N__54272\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54270\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54257\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54216\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54204\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54182\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54173\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54171\ : std_logic;
signal \N__54170\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54167\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54151\ : std_logic;
signal \N__54150\ : std_logic;
signal \N__54149\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54140\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54137\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54125\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54110\ : std_logic;
signal \N__54107\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54092\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54089\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54087\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54076\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54074\ : std_logic;
signal \N__54073\ : std_logic;
signal \N__54072\ : std_logic;
signal \N__54071\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54064\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54045\ : std_logic;
signal \N__54040\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54035\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54032\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54030\ : std_logic;
signal \N__54029\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54026\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54008\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53959\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53955\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53930\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53918\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53914\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53869\ : std_logic;
signal \N__53866\ : std_logic;
signal \N__53863\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53844\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53801\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53722\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53683\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53643\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53591\ : std_logic;
signal \N__53590\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53588\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53581\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53569\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53566\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53558\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53554\ : std_logic;
signal \N__53553\ : std_logic;
signal \N__53550\ : std_logic;
signal \N__53549\ : std_logic;
signal \N__53548\ : std_logic;
signal \N__53545\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53519\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53513\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53505\ : std_logic;
signal \N__53504\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53498\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53495\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53489\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53467\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53465\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53443\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53427\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53341\ : std_logic;
signal \N__53338\ : std_logic;
signal \N__53333\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53274\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53186\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53183\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53163\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53157\ : std_logic;
signal \N__53156\ : std_logic;
signal \N__53153\ : std_logic;
signal \N__53146\ : std_logic;
signal \N__53143\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53097\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53044\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52994\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52959\ : std_logic;
signal \N__52958\ : std_logic;
signal \N__52955\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52912\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52850\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52838\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52829\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52819\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52758\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52753\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52750\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52747\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52721\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52717\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52696\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52662\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52633\ : std_logic;
signal \N__52630\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52529\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52517\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52511\ : std_logic;
signal \N__52508\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52436\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52403\ : std_logic;
signal \N__52400\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52336\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52289\ : std_logic;
signal \N__52286\ : std_logic;
signal \N__52283\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52157\ : std_logic;
signal \N__52154\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52120\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52094\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52088\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52085\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52053\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51988\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51845\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51839\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51835\ : std_logic;
signal \N__51832\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51692\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51593\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51584\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51549\ : std_logic;
signal \N__51546\ : std_logic;
signal \N__51543\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51527\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51407\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51308\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51230\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51202\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51157\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51095\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51073\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51064\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51036\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50854\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50683\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46223\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \ADC_VAC.n19408\ : std_logic;
signal \ADC_VAC.n19409\ : std_logic;
signal \ADC_VAC.n19410\ : std_logic;
signal \ADC_VAC.n19411\ : std_logic;
signal \ADC_VAC.n19412\ : std_logic;
signal \ADC_VAC.n19413\ : std_logic;
signal \ADC_VAC.n19414\ : std_logic;
signal \ADC_VAC.bit_cnt_0\ : std_logic;
signal \ADC_VAC.bit_cnt_6\ : std_logic;
signal \ADC_VAC.bit_cnt_4\ : std_logic;
signal \ADC_VAC.bit_cnt_3\ : std_logic;
signal \ADC_VAC.bit_cnt_5\ : std_logic;
signal \ADC_VAC.bit_cnt_2\ : std_logic;
signal \ADC_VAC.bit_cnt_7\ : std_logic;
signal \ADC_VAC.bit_cnt_1\ : std_logic;
signal \ADC_VAC.n21054_cascade_\ : std_logic;
signal \ADC_VAC.n16\ : std_logic;
signal \VAC_MISO\ : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal \ADC_VAC.n14822\ : std_logic;
signal \ADC_VAC.n20715_cascade_\ : std_logic;
signal \ADC_VAC.n21053\ : std_logic;
signal \ADC_VAC.n20716\ : std_logic;
signal \ADC_VAC.n17_cascade_\ : std_logic;
signal \ADC_VAC.n12\ : std_logic;
signal \ADC_VAC.n12489\ : std_logic;
signal \VAC_SCLK\ : std_logic;
signal \n14_adj_1606_cascade_\ : std_logic;
signal \VAC_CS\ : std_logic;
signal n20615 : std_logic;
signal \VAC_DRDY\ : std_logic;
signal \n20615_cascade_\ : std_logic;
signal bit_cnt_2 : std_logic;
signal bit_cnt_1 : std_logic;
signal \CLK_DDS.n16766\ : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \ADC_VDC.n19457\ : std_logic;
signal \ADC_VDC.n19458\ : std_logic;
signal \ADC_VDC.n19459\ : std_logic;
signal \ADC_VDC.n19460\ : std_logic;
signal \ADC_VDC.n19461\ : std_logic;
signal \ADC_VDC.n19462\ : std_logic;
signal \ADC_VDC.n19463\ : std_logic;
signal \ADC_VDC.n19464\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \ADC_VDC.n19465\ : std_logic;
signal \ADC_VDC.n19466\ : std_logic;
signal \ADC_VDC.n19467\ : std_logic;
signal \ADC_VDC.avg_cnt_4\ : std_logic;
signal \ADC_VDC.avg_cnt_7\ : std_logic;
signal \ADC_VDC.avg_cnt_3\ : std_logic;
signal \ADC_VDC.avg_cnt_5\ : std_logic;
signal \ADC_VDC.avg_cnt_9\ : std_logic;
signal \ADC_VDC.avg_cnt_0\ : std_logic;
signal \ADC_VDC.avg_cnt_8\ : std_logic;
signal \ADC_VDC.avg_cnt_10\ : std_logic;
signal \ADC_VDC.n20\ : std_logic;
signal \ADC_VDC.n19_adj_1412_cascade_\ : std_logic;
signal \ADC_VDC.n18479_cascade_\ : std_logic;
signal \DDS_CS1\ : std_logic;
signal \RTD_SDO\ : std_logic;
signal \CLK_DDS.tmp_buf_0\ : std_logic;
signal bit_cnt_3 : std_logic;
signal bit_cnt_0_adj_1456 : std_logic;
signal \ADC_IAC.n17_cascade_\ : std_logic;
signal \DDS_SCK1\ : std_logic;
signal cmd_rdadctmp_6_adj_1444 : std_logic;
signal \ADC_IAC.n12\ : std_logic;
signal \n20612_cascade_\ : std_logic;
signal \ADC_IAC.n20713\ : std_logic;
signal \ADC_IAC.n20783_cascade_\ : std_logic;
signal \ADC_IAC.n20795_cascade_\ : std_logic;
signal \ADC_IAC.n21068_cascade_\ : std_logic;
signal \ADC_IAC.n20714\ : std_logic;
signal \IAC_MISO\ : std_logic;
signal cmd_rdadctmp_0_adj_1450 : std_logic;
signal \IAC_SCLK\ : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \ADC_VDC.n19531\ : std_logic;
signal \ADC_VDC.n19532\ : std_logic;
signal \ADC_VDC.n19533\ : std_logic;
signal \ADC_VDC.n19534\ : std_logic;
signal \ADC_VDC.n19535\ : std_logic;
signal \ADC_VDC.n19536\ : std_logic;
signal \ADC_VDC.n19537\ : std_logic;
signal \ADC_VDC.bit_cnt_5\ : std_logic;
signal \ADC_VDC.n20534_cascade_\ : std_logic;
signal \ADC_VDC.n10\ : std_logic;
signal \ADC_VDC.bit_cnt_7\ : std_logic;
signal \ADC_VDC.bit_cnt_6\ : std_logic;
signal \ADC_VDC.n21082\ : std_logic;
signal \ADC_VDC.n21079\ : std_logic;
signal \ADC_VDC.n21977_cascade_\ : std_logic;
signal \ADC_VDC.n18482\ : std_logic;
signal \ADC_VDC.bit_cnt_2\ : std_logic;
signal \ADC_VDC.n6\ : std_logic;
signal \ADC_VDC.n10552_cascade_\ : std_logic;
signal \ADC_VDC.n21974\ : std_logic;
signal \ADC_VDC.bit_cnt_3\ : std_logic;
signal \ADC_VDC.n20562\ : std_logic;
signal \ADC_VDC.n21224_cascade_\ : std_logic;
signal \ADC_VDC.n20748\ : std_logic;
signal \ADC_VDC.n31_cascade_\ : std_logic;
signal \ADC_VDC.n20555\ : std_logic;
signal read_buf_12 : std_logic;
signal adress_3 : std_logic;
signal adress_2 : std_logic;
signal adress_4 : std_logic;
signal adress_5 : std_logic;
signal \RTD_SDI\ : std_logic;
signal \RTD.n21309_cascade_\ : std_logic;
signal \RTD.n12\ : std_logic;
signal \RTD.n19_cascade_\ : std_logic;
signal read_buf_9 : std_logic;
signal adress_1 : std_logic;
signal read_buf_1 : std_logic;
signal read_buf_13 : std_logic;
signal read_buf_8 : std_logic;
signal n20754 : std_logic;
signal cmd_rdadctmp_5_adj_1445 : std_logic;
signal cmd_rdadctmp_4_adj_1446 : std_logic;
signal cmd_rdadctmp_3_adj_1447 : std_logic;
signal \IAC_DRDY\ : std_logic;
signal n20612 : std_logic;
signal \n14_adj_1604_cascade_\ : std_logic;
signal \IAC_CS\ : std_logic;
signal \ADC_IAC.bit_cnt_0\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \ADC_IAC.bit_cnt_1\ : std_logic;
signal \ADC_IAC.n19415\ : std_logic;
signal \ADC_IAC.bit_cnt_2\ : std_logic;
signal \ADC_IAC.n19416\ : std_logic;
signal \ADC_IAC.bit_cnt_3\ : std_logic;
signal \ADC_IAC.n19417\ : std_logic;
signal \ADC_IAC.bit_cnt_4\ : std_logic;
signal \ADC_IAC.n19418\ : std_logic;
signal \ADC_IAC.bit_cnt_5\ : std_logic;
signal \ADC_IAC.n19419\ : std_logic;
signal \ADC_IAC.bit_cnt_6\ : std_logic;
signal \ADC_IAC.n19420\ : std_logic;
signal \ADC_IAC.n19421\ : std_logic;
signal \ADC_IAC.bit_cnt_7\ : std_logic;
signal \ADC_IAC.n12586\ : std_logic;
signal \ADC_IAC.n14860\ : std_logic;
signal cmd_rdadctmp_1_adj_1449 : std_logic;
signal cmd_rdadctmp_2_adj_1448 : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal cmd_rdadctmp_28_adj_1422 : std_logic;
signal \ADC_VDC.n19_adj_1413_cascade_\ : std_logic;
signal \ADC_VDC.n17\ : std_logic;
signal \ADC_VDC.n4\ : std_logic;
signal \ADC_VDC.n10132_cascade_\ : std_logic;
signal \ADC_VDC.n7_adj_1411\ : std_logic;
signal \ADC_VDC.n20750\ : std_logic;
signal \ADC_VDC.n12\ : std_logic;
signal \ADC_VDC.n20750_cascade_\ : std_logic;
signal \ADC_VDC.n11692_cascade_\ : std_logic;
signal \VDC_SCLK\ : std_logic;
signal \ADC_VDC.bit_cnt_1\ : std_logic;
signal \ADC_VDC.n20534\ : std_logic;
signal \ADC_VDC.bit_cnt_4\ : std_logic;
signal \ADC_VDC.n6_adj_1410\ : std_logic;
signal \ADC_VDC.n11281_cascade_\ : std_logic;
signal \ADC_VDC.bit_cnt_0\ : std_logic;
signal \ADC_VDC.n15\ : std_logic;
signal \ADC_VDC.n15_cascade_\ : std_logic;
signal \ADC_VDC.n20746_cascade_\ : std_logic;
signal \ADC_VDC.n72\ : std_logic;
signal \ADC_VDC.n12823\ : std_logic;
signal \ADC_VDC.n13038_cascade_\ : std_logic;
signal \ADC_VDC.n20659\ : std_logic;
signal \ADC_VDC.n17432_cascade_\ : std_logic;
signal \ADC_VDC.n18466\ : std_logic;
signal read_buf_11 : std_logic;
signal read_buf_15 : std_logic;
signal \n11730_cascade_\ : std_logic;
signal adress_6 : std_logic;
signal \RTD.cfg_buf_6\ : std_logic;
signal \RTD.cfg_buf_0\ : std_logic;
signal \RTD.n9_cascade_\ : std_logic;
signal \RTD.adress_7_N_1340_7_cascade_\ : std_logic;
signal \RTD.adress_7\ : std_logic;
signal adress_0 : std_logic;
signal n13181 : std_logic;
signal \RTD.cfg_buf_5\ : std_logic;
signal \RTD.cfg_buf_3\ : std_logic;
signal \RTD.n11\ : std_logic;
signal \RTD.n7333_cascade_\ : std_logic;
signal \RTD.n13_cascade_\ : std_logic;
signal \RTD.n11734\ : std_logic;
signal \RTD.n7333\ : std_logic;
signal \RTD.cfg_tmp_1\ : std_logic;
signal \RTD.cfg_tmp_2\ : std_logic;
signal \RTD.cfg_tmp_3\ : std_logic;
signal \RTD.cfg_tmp_4\ : std_logic;
signal \RTD.cfg_tmp_5\ : std_logic;
signal \RTD.cfg_tmp_6\ : std_logic;
signal \RTD.cfg_tmp_7\ : std_logic;
signal \RTD.cfg_tmp_0\ : std_logic;
signal \RTD.n13228\ : std_logic;
signal \RTD.n15015\ : std_logic;
signal read_buf_7 : std_logic;
signal read_buf_2 : std_logic;
signal read_buf_3 : std_logic;
signal n1_adj_1601 : std_logic;
signal read_buf_4 : std_logic;
signal \n1_adj_1601_cascade_\ : std_logic;
signal read_buf_5 : std_logic;
signal cmd_rdadctmp_29_adj_1421 : std_logic;
signal cmd_rdadctmp_30_adj_1420 : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal cmd_rdadctmp_23_adj_1427 : std_logic;
signal cmd_rdadctmp_24_adj_1426 : std_logic;
signal cmd_rdadctmp_26_adj_1424 : std_logic;
signal \CLK_DDS.tmp_buf_1\ : std_logic;
signal \CLK_DDS.tmp_buf_2\ : std_logic;
signal \CLK_DDS.tmp_buf_3\ : std_logic;
signal \CLK_DDS.tmp_buf_4\ : std_logic;
signal \CLK_DDS.tmp_buf_5\ : std_logic;
signal \CLK_DDS.tmp_buf_6\ : std_logic;
signal \CLK_DDS.tmp_buf_7\ : std_logic;
signal \CLK_DDS.n9_adj_1395\ : std_logic;
signal buf_adcdata_vac_4 : std_logic;
signal \n19_adj_1636_cascade_\ : std_logic;
signal buf_adcdata_iac_4 : std_logic;
signal buf_data_iac_4 : std_logic;
signal \n22_adj_1637_cascade_\ : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal n19_adj_1631 : std_logic;
signal buf_adcdata_vac_5 : std_logic;
signal buf_adcdata_vac_20 : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal buf_adcdata_vdc_5 : std_logic;
signal buf_adcdata_vdc_4 : std_logic;
signal buf_adcdata_vdc_20 : std_logic;
signal \ADC_VDC.n47\ : std_logic;
signal \RTD_SCLK\ : std_logic;
signal \RTD.n8\ : std_logic;
signal n13309 : std_logic;
signal \RTD_DRDY\ : std_logic;
signal \RTD.adress_7_N_1340_7\ : std_logic;
signal \RTD.n16669\ : std_logic;
signal \RTD.n16669_cascade_\ : std_logic;
signal \RTD_CS\ : std_logic;
signal \RTD.n11703\ : std_logic;
signal \RTD.cfg_buf_1\ : std_logic;
signal \RTD.n12_adj_1397\ : std_logic;
signal buf_adcdata_vdc_23 : std_logic;
signal buf_adcdata_vac_23 : std_logic;
signal \n19_adj_1526_cascade_\ : std_logic;
signal \n22076_cascade_\ : std_logic;
signal \buf_readRTD_15\ : std_logic;
signal n20 : std_logic;
signal \RTD.n22370\ : std_logic;
signal \RTD.n21323_cascade_\ : std_logic;
signal \RTD.n26\ : std_logic;
signal \RTD.n21325_cascade_\ : std_logic;
signal \RTD.n4\ : std_logic;
signal \RTD.n1\ : std_logic;
signal \RTD.n1_cascade_\ : std_logic;
signal \RTD.n20587\ : std_logic;
signal n8_adj_1608 : std_logic;
signal n21227 : std_logic;
signal dds_state_0_adj_1454 : std_logic;
signal \CLK_DDS.n9\ : std_logic;
signal \RTD.mode\ : std_logic;
signal \RTD.n21276_cascade_\ : std_logic;
signal \RTD.n21275\ : std_logic;
signal \RTD.adc_state_3_N_1368_1\ : std_logic;
signal \RTD.adc_state_3_N_1368_1_cascade_\ : std_logic;
signal \RTD.n7\ : std_logic;
signal \RTD.n20762\ : std_logic;
signal \RTD.n11742\ : std_logic;
signal \n16_adj_1512_cascade_\ : std_logic;
signal cmd_rdadctmp_25_adj_1425 : std_logic;
signal cmd_rdadctmp_31_adj_1419 : std_logic;
signal \VAC_OSR1\ : std_logic;
signal buf_adcdata_iac_21 : std_logic;
signal buf_adcdata_iac_23 : std_logic;
signal \VAC_FLT1\ : std_logic;
signal n17_adj_1525 : std_logic;
signal buf_adcdata_iac_16 : std_logic;
signal \IAC_OSR0\ : std_logic;
signal n22100 : std_logic;
signal \SELIRNG0\ : std_logic;
signal \CLK_DDS.tmp_buf_10\ : std_logic;
signal \CLK_DDS.tmp_buf_11\ : std_logic;
signal \CLK_DDS.tmp_buf_12\ : std_logic;
signal \CLK_DDS.tmp_buf_13\ : std_logic;
signal \CLK_DDS.tmp_buf_14\ : std_logic;
signal tmp_buf_15_adj_1455 : std_logic;
signal dds_state_2_adj_1452 : std_logic;
signal dds_state_1_adj_1453 : std_logic;
signal \CLK_DDS.tmp_buf_8\ : std_logic;
signal \CLK_DDS.tmp_buf_9\ : std_logic;
signal \CLK_DDS.n12800\ : std_logic;
signal trig_dds1 : std_logic;
signal \ICE_GPMO_1\ : std_logic;
signal \IAC_CLK\ : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal buf_adcdata_vdc_7 : std_logic;
signal buf_adcdata_vac_7 : std_logic;
signal buf_adcdata_iac_7 : std_logic;
signal \n19_adj_1625_cascade_\ : std_logic;
signal buf_data_iac_7 : std_logic;
signal \n22_adj_1626_cascade_\ : std_logic;
signal buf_adcdata_vac_6 : std_logic;
signal buf_adcdata_vdc_6 : std_logic;
signal buf_adcdata_iac_6 : std_logic;
signal \n19_adj_1628_cascade_\ : std_logic;
signal buf_data_iac_6 : std_logic;
signal \n22_adj_1629_cascade_\ : std_logic;
signal cmd_rdadctmp_14_adj_1436 : std_logic;
signal cmd_rdadctmp_15_adj_1435 : std_logic;
signal \n12875_cascade_\ : std_logic;
signal buf_adcdata_vdc_19 : std_logic;
signal \ADC_VDC.avg_cnt_11\ : std_logic;
signal \ADC_VDC.avg_cnt_2\ : std_logic;
signal \ADC_VDC.avg_cnt_1\ : std_logic;
signal \ADC_VDC.avg_cnt_6\ : std_logic;
signal \ADC_VDC.n21\ : std_logic;
signal \ADC_VDC.n18479\ : std_logic;
signal \ADC_VDC.n21145_cascade_\ : std_logic;
signal \ADC_VDC.n13050\ : std_logic;
signal read_buf_10 : std_logic;
signal buf_adcdata_vdc_18 : std_logic;
signal \n20833_cascade_\ : std_logic;
signal read_buf_14 : std_logic;
signal \buf_readRTD_11\ : std_logic;
signal n22214 : std_logic;
signal \RTD.n10\ : std_logic;
signal \RTD.cfg_buf_2\ : std_logic;
signal read_buf_0 : std_logic;
signal \RTD.adc_state_0\ : std_logic;
signal adc_state_3_adj_1481 : std_logic;
signal \RTD.n14717\ : std_logic;
signal n16_adj_1524 : std_logic;
signal \RTD.cfg_buf_4\ : std_logic;
signal adc_state_2_adj_1482 : std_logic;
signal read_buf_6 : std_logic;
signal n11730 : std_logic;
signal \RTD.n13192\ : std_logic;
signal \RTD.n20631\ : std_logic;
signal \buf_cfgRTD_7\ : std_logic;
signal \RTD.cfg_buf_7\ : std_logic;
signal \buf_cfgRTD_3\ : std_logic;
signal cmd_rdadctmp_7_adj_1443 : std_logic;
signal \buf_readRTD_13\ : std_logic;
signal \buf_readRTD_10\ : std_logic;
signal \buf_cfgRTD_2\ : std_logic;
signal n20834 : std_logic;
signal adc_state_1_adj_1483 : std_logic;
signal \RTD.n20656\ : std_logic;
signal \n12397_cascade_\ : std_logic;
signal buf_adcdata_vac_21 : std_logic;
signal buf_adcdata_vdc_21 : std_logic;
signal n22184 : std_logic;
signal \buf_readRTD_12\ : std_logic;
signal n22202 : std_logic;
signal \buf_readRTD_8\ : std_logic;
signal \buf_cfgRTD_0\ : std_logic;
signal cmd_rdadctmp_27_adj_1423 : std_logic;
signal buf_dds1_15 : std_logic;
signal \buf_cfgRTD_4\ : std_logic;
signal n20849 : std_logic;
signal n22103 : std_logic;
signal buf_adcdata_iac_17 : std_logic;
signal buf_data_iac_21 : std_logic;
signal \n20876_cascade_\ : std_logic;
signal n22106 : std_logic;
signal n20875 : std_logic;
signal n22022 : std_logic;
signal buf_dds1_4 : std_logic;
signal \n8_adj_1555_cascade_\ : std_logic;
signal \data_index_9_N_216_8\ : std_logic;
signal n8_adj_1555 : std_logic;
signal n22040 : std_logic;
signal buf_dds1_9 : std_logic;
signal buf_dds1_8 : std_logic;
signal \n12383_cascade_\ : std_logic;
signal buf_dds1_10 : std_logic;
signal n20673 : std_logic;
signal \n11412_cascade_\ : std_logic;
signal \AC_ADC_SYNC\ : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal cmd_rdadctmp_13_adj_1437 : std_logic;
signal buf_adcdata_iac_5 : std_logic;
signal buf_data_iac_5 : std_logic;
signal n22_adj_1632 : std_logic;
signal \ADC_VDC.n21718\ : std_logic;
signal n12875 : std_logic;
signal cmd_rdadctmp_0_adj_1479 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_0\ : std_logic;
signal \bfn_10_5_0_\ : std_logic;
signal cmd_rdadctmp_1_adj_1478 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_1\ : std_logic;
signal \ADC_VDC.n19422\ : std_logic;
signal cmd_rdadctmp_2_adj_1477 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_2\ : std_logic;
signal \ADC_VDC.n19423\ : std_logic;
signal cmd_rdadctmp_3_adj_1476 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_3\ : std_logic;
signal \ADC_VDC.n19424\ : std_logic;
signal cmd_rdadctmp_4_adj_1475 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_4\ : std_logic;
signal \ADC_VDC.n19425\ : std_logic;
signal cmd_rdadctmp_5_adj_1474 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_5\ : std_logic;
signal \ADC_VDC.n19426\ : std_logic;
signal cmd_rdadctmp_6_adj_1473 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_6\ : std_logic;
signal \ADC_VDC.n19427\ : std_logic;
signal cmd_rdadctmp_7_adj_1472 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_7\ : std_logic;
signal \ADC_VDC.n19428\ : std_logic;
signal \ADC_VDC.n19429\ : std_logic;
signal cmd_rdadctmp_8_adj_1471 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_8\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal cmd_rdadctmp_9_adj_1470 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_9\ : std_logic;
signal \ADC_VDC.n19430\ : std_logic;
signal cmd_rdadctmp_10_adj_1469 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_10\ : std_logic;
signal \ADC_VDC.n19431\ : std_logic;
signal cmd_rdadctmp_11_adj_1468 : std_logic;
signal \ADC_VDC.n19432\ : std_logic;
signal cmd_rdadctmp_12_adj_1467 : std_logic;
signal cmd_rdadcbuf_12 : std_logic;
signal \ADC_VDC.n19433\ : std_logic;
signal cmd_rdadctmp_13_adj_1466 : std_logic;
signal cmd_rdadcbuf_13 : std_logic;
signal \ADC_VDC.n19434\ : std_logic;
signal cmd_rdadctmp_14_adj_1465 : std_logic;
signal cmd_rdadcbuf_14 : std_logic;
signal \ADC_VDC.n19435\ : std_logic;
signal cmd_rdadctmp_15_adj_1464 : std_logic;
signal cmd_rdadcbuf_15 : std_logic;
signal \ADC_VDC.n19436\ : std_logic;
signal \ADC_VDC.n19437\ : std_logic;
signal cmd_rdadctmp_16_adj_1463 : std_logic;
signal cmd_rdadcbuf_16 : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal cmd_rdadctmp_17_adj_1462 : std_logic;
signal cmd_rdadcbuf_17 : std_logic;
signal \ADC_VDC.n19438\ : std_logic;
signal cmd_rdadctmp_18_adj_1461 : std_logic;
signal cmd_rdadcbuf_18 : std_logic;
signal \ADC_VDC.n19439\ : std_logic;
signal cmd_rdadctmp_19_adj_1460 : std_logic;
signal cmd_rdadcbuf_19 : std_logic;
signal \ADC_VDC.n19440\ : std_logic;
signal cmd_rdadctmp_20_adj_1459 : std_logic;
signal \ADC_VDC.n19441\ : std_logic;
signal cmd_rdadctmp_21_adj_1458 : std_logic;
signal cmd_rdadcbuf_21 : std_logic;
signal \ADC_VDC.n19442\ : std_logic;
signal cmd_rdadcbuf_22 : std_logic;
signal \ADC_VDC.n19443\ : std_logic;
signal cmd_rdadcbuf_23 : std_logic;
signal \ADC_VDC.n19444\ : std_logic;
signal \ADC_VDC.n19445\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \ADC_VDC.n19446\ : std_logic;
signal \ADC_VDC.n19447\ : std_logic;
signal \ADC_VDC.n19448\ : std_logic;
signal cmd_rdadcbuf_28 : std_logic;
signal \ADC_VDC.n19449\ : std_logic;
signal cmd_rdadcbuf_29 : std_logic;
signal \ADC_VDC.n19450\ : std_logic;
signal cmd_rdadcbuf_30 : std_logic;
signal \ADC_VDC.n19451\ : std_logic;
signal cmd_rdadcbuf_31 : std_logic;
signal \ADC_VDC.n19452\ : std_logic;
signal \ADC_VDC.n19453\ : std_logic;
signal cmd_rdadcbuf_32 : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \ADC_VDC.n19454\ : std_logic;
signal \ADC_VDC.n13038\ : std_logic;
signal \ADC_VDC.n14931\ : std_logic;
signal cmd_rdadcbuf_34 : std_logic;
signal \ADC_VDC.n19455\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_35_N_1139_34\ : std_logic;
signal n20824 : std_logic;
signal n22118 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal \buf_cfgRTD_5\ : std_logic;
signal buf_adcdata_iac_18 : std_logic;
signal \IAC_FLT0\ : std_logic;
signal n20825 : std_logic;
signal \data_index_9_N_216_0\ : std_logic;
signal comm_cmd_5 : std_logic;
signal comm_cmd_6 : std_logic;
signal \IAC_OSR1\ : std_logic;
signal comm_cmd_4 : std_logic;
signal buf_dds1_3 : std_logic;
signal \buf_cfgRTD_1\ : std_logic;
signal \buf_readRTD_9\ : std_logic;
signal n9_adj_1416 : std_logic;
signal buf_dds1_0 : std_logic;
signal \n20663_cascade_\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal n19384 : std_logic;
signal n19385 : std_logic;
signal n19386 : std_logic;
signal n19387 : std_logic;
signal n19388 : std_logic;
signal n19389 : std_logic;
signal n19390 : std_logic;
signal n19391 : std_logic;
signal data_index_8 : std_logic;
signal n7_adj_1554 : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal n19392 : std_logic;
signal buf_dds1_2 : std_logic;
signal data_index_7 : std_logic;
signal n8_adj_1557 : std_logic;
signal \n8_adj_1557_cascade_\ : std_logic;
signal n7_adj_1556 : std_logic;
signal \data_index_9_N_216_7\ : std_logic;
signal \n8_adj_1553_cascade_\ : std_logic;
signal data_index_9 : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal n11401 : std_logic;
signal \n20772_cascade_\ : std_logic;
signal \n11835_cascade_\ : std_logic;
signal buf_dds0_10 : std_logic;
signal \SIG_DDS.tmp_buf_10\ : std_logic;
signal buf_dds0_13 : std_logic;
signal \SIG_DDS.tmp_buf_13\ : std_logic;
signal \SIG_DDS.tmp_buf_11\ : std_logic;
signal \SIG_DDS.tmp_buf_12\ : std_logic;
signal \SIG_DDS.tmp_buf_14\ : std_logic;
signal buf_dds0_15 : std_logic;
signal buf_dds0_9 : std_logic;
signal \SIG_DDS.tmp_buf_9\ : std_logic;
signal \SIG_DDS.tmp_buf_6\ : std_logic;
signal \SIG_DDS.tmp_buf_5\ : std_logic;
signal buf_dds0_2 : std_logic;
signal buf_dds0_4 : std_logic;
signal \SIG_DDS.tmp_buf_4\ : std_logic;
signal \SIG_DDS.tmp_buf_7\ : std_logic;
signal buf_dds0_8 : std_logic;
signal \SIG_DDS.tmp_buf_8\ : std_logic;
signal buf_dds0_1 : std_logic;
signal \SIG_DDS.tmp_buf_1\ : std_logic;
signal \SIG_DDS.tmp_buf_2\ : std_logic;
signal buf_dds0_3 : std_logic;
signal \SIG_DDS.tmp_buf_3\ : std_logic;
signal n8_adj_1553 : std_logic;
signal n7_adj_1552 : std_logic;
signal \data_index_9_N_216_9\ : std_logic;
signal buf_adcdata_vdc_2 : std_logic;
signal buf_adcdata_vac_2 : std_logic;
signal buf_adcdata_iac_2 : std_logic;
signal \n19_adj_1646_cascade_\ : std_logic;
signal buf_data_iac_2 : std_logic;
signal \n22_adj_1647_cascade_\ : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal buf_adcdata_vdc_3 : std_logic;
signal \n19_adj_1642_cascade_\ : std_logic;
signal buf_data_iac_3 : std_logic;
signal \n22_adj_1643_cascade_\ : std_logic;
signal buf_adcdata_iac_3 : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal buf_adcdata_vac_3 : std_logic;
signal cmd_rdadctmp_11_adj_1439 : std_logic;
signal cmd_rdadctmp_12_adj_1438 : std_logic;
signal buf_data_vac_7 : std_logic;
signal buf_data_vac_6 : std_logic;
signal buf_data_vac_5 : std_logic;
signal cmd_rdadctmp_10_adj_1440 : std_logic;
signal \n30_adj_1480_cascade_\ : std_logic;
signal buf_adcdata_vdc_1 : std_logic;
signal \n19_adj_1491_cascade_\ : std_logic;
signal buf_adcdata_iac_1 : std_logic;
signal \buf_readRTD_14\ : std_logic;
signal cmd_rdadcbuf_26 : std_logic;
signal cmd_rdadcbuf_25 : std_logic;
signal cmd_rdadcbuf_24 : std_logic;
signal cmd_rdadcbuf_27 : std_logic;
signal cmd_rdadcbuf_11 : std_logic;
signal cmd_rdadcbuf_33 : std_logic;
signal n13109 : std_logic;
signal cmd_rdadcbuf_20 : std_logic;
signal buf_adcdata_vac_18 : std_logic;
signal n12411 : std_logic;
signal \buf_cfgRTD_6\ : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal buf_adcdata_vac_19 : std_logic;
signal cmd_rdadctmp_8_adj_1442 : std_logic;
signal cmd_rdadctmp_9_adj_1441 : std_logic;
signal buf_adcdata_vdc_15 : std_logic;
signal buf_adcdata_vac_15 : std_logic;
signal n22016 : std_logic;
signal buf_adcdata_vdc_16 : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal \n20590_cascade_\ : std_logic;
signal buf_adcdata_vac_16 : std_logic;
signal data_count_0 : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n19345 : std_logic;
signal data_count_2 : std_logic;
signal n19346 : std_logic;
signal data_count_3 : std_logic;
signal n19347 : std_logic;
signal data_count_4 : std_logic;
signal n19348 : std_logic;
signal data_count_5 : std_logic;
signal n19349 : std_logic;
signal data_count_6 : std_logic;
signal n19350 : std_logic;
signal data_count_7 : std_logic;
signal n19351 : std_logic;
signal n19352 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal data_count_8 : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal n19353 : std_logic;
signal data_count_9 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal buf_adcdata_vdc_8 : std_logic;
signal buf_adcdata_vac_8 : std_logic;
signal buf_adcdata_vdc_10 : std_logic;
signal buf_adcdata_vac_10 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal \AMPV_POW\ : std_logic;
signal n23_adj_1536 : std_logic;
signal cmd_rdadctmp_21_adj_1429 : std_logic;
signal n7_adj_1531 : std_logic;
signal cmd_rdadctmp_22_adj_1428 : std_logic;
signal buf_adcdata_vdc_9 : std_logic;
signal buf_adcdata_vac_9 : std_logic;
signal \n17411_cascade_\ : std_logic;
signal \data_index_9_N_216_5\ : std_logic;
signal n17409 : std_logic;
signal n17411 : std_logic;
signal data_index_5 : std_logic;
signal \n8828_cascade_\ : std_logic;
signal data_index_0 : std_logic;
signal n8_adj_1532 : std_logic;
signal buf_dds1_13 : std_logic;
signal buf_dds0_6 : std_logic;
signal buf_dds1_6 : std_logic;
signal n11757 : std_logic;
signal wdtick_cnt_0 : std_logic;
signal wdtick_cnt_1 : std_logic;
signal wdtick_cnt_2 : std_logic;
signal buf_dds0_0 : std_logic;
signal \SIG_DDS.tmp_buf_0\ : std_logic;
signal \SIG_DDS.n12738\ : std_logic;
signal \EIS_SYNCCLK\ : std_logic;
signal \OUT_SYNCCLK\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \ADC_VDC.genclk.n19468\ : std_logic;
signal \ADC_VDC.genclk.t0off_2\ : std_logic;
signal \ADC_VDC.genclk.n19469\ : std_logic;
signal \ADC_VDC.genclk.n19470\ : std_logic;
signal \ADC_VDC.genclk.n19471\ : std_logic;
signal \ADC_VDC.genclk.n19472\ : std_logic;
signal \ADC_VDC.genclk.n19473\ : std_logic;
signal \ADC_VDC.genclk.t0off_7\ : std_logic;
signal \ADC_VDC.genclk.n19474\ : std_logic;
signal \ADC_VDC.genclk.n19475\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i0C_net\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \ADC_VDC.genclk.n19476\ : std_logic;
signal \ADC_VDC.genclk.t0off_10\ : std_logic;
signal \ADC_VDC.genclk.n19477\ : std_logic;
signal \ADC_VDC.genclk.n19478\ : std_logic;
signal \ADC_VDC.genclk.t0off_12\ : std_logic;
signal \ADC_VDC.genclk.n19479\ : std_logic;
signal \ADC_VDC.genclk.n19480\ : std_logic;
signal \ADC_VDC.genclk.n19481\ : std_logic;
signal \ADC_VDC.genclk.n19482\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.n11751\ : std_logic;
signal \n12_adj_1615_cascade_\ : std_logic;
signal \n12236_cascade_\ : std_logic;
signal buf_data_vac_0 : std_logic;
signal buf_data_vac_1 : std_logic;
signal buf_data_vac_2 : std_logic;
signal buf_data_vac_3 : std_logic;
signal buf_data_vac_4 : std_logic;
signal n12236 : std_logic;
signal n14801 : std_logic;
signal \n2_adj_1587_cascade_\ : std_logic;
signal comm_buf_5_4 : std_logic;
signal n21324 : std_logic;
signal \n4_adj_1588_cascade_\ : std_logic;
signal n22136 : std_logic;
signal n1_adj_1586 : std_logic;
signal n19006 : std_logic;
signal \n19006_cascade_\ : std_logic;
signal n30_adj_1627 : std_logic;
signal n30_adj_1630 : std_logic;
signal n30_adj_1634 : std_logic;
signal n30_adj_1638 : std_logic;
signal comm_buf_2_4 : std_logic;
signal n30_adj_1644 : std_logic;
signal n30_adj_1648 : std_logic;
signal cmd_rdadctmp_22_adj_1457 : std_logic;
signal \ADC_VDC.n10552\ : std_logic;
signal \ADC_VDC.cmd_rdadctmp_23\ : std_logic;
signal \ADC_VDC.n12915\ : std_logic;
signal \ADC_VDC.n20392\ : std_logic;
signal \RTD.n17720\ : std_logic;
signal buf_adcdata_vac_22 : std_logic;
signal buf_adcdata_vdc_22 : std_logic;
signal n22160 : std_logic;
signal comm_buf_6_4 : std_logic;
signal n20646 : std_logic;
signal n14522 : std_logic;
signal n11918 : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal n19393 : std_logic;
signal n19394 : std_logic;
signal n19395 : std_logic;
signal n19396 : std_logic;
signal n19397 : std_logic;
signal n19398 : std_logic;
signal n19399 : std_logic;
signal n19400 : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal n19401 : std_logic;
signal n19402 : std_logic;
signal n19403 : std_logic;
signal n19404 : std_logic;
signal data_idxvec_13 : std_logic;
signal n19405 : std_logic;
signal n19406 : std_logic;
signal n19407 : std_logic;
signal \n22169_cascade_\ : std_logic;
signal n22079 : std_logic;
signal \n20568_cascade_\ : std_logic;
signal data_idxvec_15 : std_logic;
signal eis_end : std_logic;
signal \n26_adj_1528_cascade_\ : std_logic;
signal n22166 : std_logic;
signal n20742 : std_logic;
signal acadc_trig : std_logic;
signal \INVeis_end_309C_net\ : std_logic;
signal \n16594_cascade_\ : std_logic;
signal n22196 : std_logic;
signal \n16602_cascade_\ : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal n16602 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n19369 : std_logic;
signal \n19369_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n19369_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n19369_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n19369_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n19369_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n19369_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n19369_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal n19370 : std_logic;
signal n19371 : std_logic;
signal n19372 : std_logic;
signal n19373 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal n19374 : std_logic;
signal n19375 : std_logic;
signal n19376 : std_logic;
signal n19377 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal n19378 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal n19379 : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal n19380 : std_logic;
signal n19381 : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal n19382 : std_logic;
signal n19383 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal \TEST_LED\ : std_logic;
signal \ADC_VDC.genclk.t0off_13\ : std_logic;
signal \ADC_VDC.genclk.t0off_3\ : std_logic;
signal \ADC_VDC.genclk.t0off_5\ : std_logic;
signal \ADC_VDC.genclk.t0off_8\ : std_logic;
signal \ADC_VDC.genclk.n27\ : std_logic;
signal \ADC_VDC.genclk.n26_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21206_cascade_\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.t0off_6\ : std_logic;
signal \ADC_VDC.genclk.t0off_0\ : std_logic;
signal \ADC_VDC.genclk.t0off_4\ : std_logic;
signal \ADC_VDC.genclk.t0off_1\ : std_logic;
signal \ADC_VDC.genclk.n21208\ : std_logic;
signal \ADC_VDC.genclk.t0off_14\ : std_logic;
signal \ADC_VDC.genclk.t0off_9\ : std_logic;
signal \ADC_VDC.genclk.t0off_15\ : std_logic;
signal \ADC_VDC.genclk.t0off_11\ : std_logic;
signal \ADC_VDC.genclk.n28\ : std_logic;
signal \ADC_VDC.genclk.n21206\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i1C_net\ : std_logic;
signal \ADC_VDC.genclk.n6\ : std_logic;
signal \ADC_VDC.genclk.div_state_0\ : std_logic;
signal \ADC_VDC.n11766\ : std_logic;
signal \VDC_SDO\ : std_logic;
signal \ADC_VDC.adc_state_0\ : std_logic;
signal \ADC_VDC.n62\ : std_logic;
signal adc_state_2 : std_logic;
signal adc_state_3 : std_logic;
signal \ADC_VDC.n62_cascade_\ : std_logic;
signal \ADC_VDC.adc_state_1\ : std_logic;
signal \ADC_VDC.n11\ : std_logic;
signal \bfn_13_5_0_\ : std_logic;
signal \ADC_VDC.genclk.n19483\ : std_logic;
signal \ADC_VDC.genclk.n19484\ : std_logic;
signal \ADC_VDC.genclk.n19485\ : std_logic;
signal \ADC_VDC.genclk.n19486\ : std_logic;
signal \ADC_VDC.genclk.n19487\ : std_logic;
signal \ADC_VDC.genclk.n19488\ : std_logic;
signal \ADC_VDC.genclk.n19489\ : std_logic;
signal \ADC_VDC.genclk.n19490\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i0C_net\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \ADC_VDC.genclk.n19491\ : std_logic;
signal \ADC_VDC.genclk.n19492\ : std_logic;
signal \ADC_VDC.genclk.n19493\ : std_logic;
signal \ADC_VDC.genclk.n19494\ : std_logic;
signal \ADC_VDC.genclk.n19495\ : std_logic;
signal \ADC_VDC.genclk.n19496\ : std_logic;
signal \ADC_VDC.genclk.n19497\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.div_state_1__N_1275\ : std_logic;
signal \ADC_VDC.genclk.n15067\ : std_logic;
signal \RTD.bit_cnt_3\ : std_logic;
signal \RTD.bit_cnt_1\ : std_logic;
signal \RTD.bit_cnt_2\ : std_logic;
signal \RTD.bit_cnt_0\ : std_logic;
signal \RTD.n11756\ : std_logic;
signal \RTD.n15081\ : std_logic;
signal \n12152_cascade_\ : std_logic;
signal n12_adj_1639 : std_logic;
signal \n12194_cascade_\ : std_logic;
signal buf_adcdata_iac_0 : std_logic;
signal \n22_cascade_\ : std_logic;
signal buf_data_iac_0 : std_logic;
signal \n30_adj_1484_cascade_\ : std_logic;
signal n22_adj_1489 : std_logic;
signal buf_data_iac_1 : std_logic;
signal \n30_adj_1504_cascade_\ : std_logic;
signal buf_adcdata_vdc_0 : std_logic;
signal buf_adcdata_vac_0 : std_logic;
signal n19_adj_1485 : std_logic;
signal n12110 : std_logic;
signal \n12110_cascade_\ : std_logic;
signal n14780 : std_logic;
signal data_idxvec_10 : std_logic;
signal \n20905_cascade_\ : std_logic;
signal n20839 : std_logic;
signal \n22148_cascade_\ : std_logic;
signal n22121 : std_logic;
signal \n22151_cascade_\ : std_logic;
signal \n20889_cascade_\ : std_logic;
signal buf_data_iac_18 : std_logic;
signal n20906 : std_logic;
signal n20670 : std_logic;
signal n20672 : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal buf_adcdata_vac_1 : std_logic;
signal n20840 : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal n20590 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal n12534 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal \n24_adj_1622_cascade_\ : std_logic;
signal buf_adcdata_vdc_12 : std_logic;
signal buf_adcdata_vac_12 : std_logic;
signal \n35_cascade_\ : std_logic;
signal \iac_raw_buf_N_735\ : std_logic;
signal n17_adj_1645 : std_logic;
signal adc_state_0 : std_logic;
signal adc_state_1 : std_logic;
signal \DTRIG_N_919\ : std_logic;
signal n8 : std_logic;
signal n11354 : std_logic;
signal \n10534_cascade_\ : std_logic;
signal n16598 : std_logic;
signal n20957 : std_logic;
signal \DTRIG_N_919_adj_1451\ : std_logic;
signal adc_state_1_adj_1417 : std_logic;
signal \ICE_GPMO_0\ : std_logic;
signal auxmode : std_logic;
signal \acadc_rst_cascade_\ : std_logic;
signal tacadc_rst : std_logic;
signal \buf_readRTD_7\ : std_logic;
signal n19_adj_1502 : std_logic;
signal \n11_cascade_\ : std_logic;
signal \n21099_cascade_\ : std_logic;
signal n13 : std_logic;
signal \INVeis_state_i2C_net\ : std_logic;
signal n11760 : std_logic;
signal n17430 : std_logic;
signal acadc_dtrig_v : std_logic;
signal acadc_dtrig_i : std_logic;
signal n4_adj_1569 : std_logic;
signal data_index_3 : std_logic;
signal n8_adj_1563 : std_logic;
signal \n8_adj_1563_cascade_\ : std_logic;
signal n7_adj_1562 : std_logic;
signal \data_index_9_N_216_3\ : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal \n20_adj_1617_cascade_\ : std_logic;
signal n17_adj_1612 : std_logic;
signal \n26_adj_1640_cascade_\ : std_logic;
signal n31 : std_logic;
signal data_index_2 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal n21 : std_logic;
signal \n24_adj_1537_cascade_\ : std_logic;
signal n23_adj_1624 : std_logic;
signal n30 : std_logic;
signal n20789 : std_logic;
signal eis_state_0 : std_logic;
signal acadc_rst : std_logic;
signal buf_dds1_5 : std_logic;
signal data_idxvec_14 : std_logic;
signal \eis_end_N_725\ : std_logic;
signal n11670 : std_logic;
signal n14687 : std_logic;
signal n10733 : std_logic;
signal buf_dds0_5 : std_logic;
signal \n27_adj_1551_cascade_\ : std_logic;
signal n25 : std_logic;
signal \n19608_cascade_\ : std_logic;
signal n10_adj_1594 : std_logic;
signal n26_adj_1543 : std_logic;
signal n28_adj_1621 : std_logic;
signal n14_adj_1592 : std_logic;
signal buf_dds1_14 : std_logic;
signal buf_dds0_14 : std_logic;
signal \n22115_cascade_\ : std_logic;
signal n22163 : std_logic;
signal \VAC_FLT0\ : std_logic;
signal buf_adcdata_iac_22 : std_logic;
signal n22112 : std_logic;
signal n21037 : std_logic;
signal n23_adj_1534 : std_logic;
signal \n22070_cascade_\ : std_logic;
signal n20856 : std_logic;
signal \n22073_cascade_\ : std_logic;
signal \n30_adj_1535_cascade_\ : std_logic;
signal \ADC_VDC.genclk.t0on_6\ : std_logic;
signal \ADC_VDC.genclk.t0on_1\ : std_logic;
signal \ADC_VDC.genclk.t0on_4\ : std_logic;
signal \ADC_VDC.genclk.t0on_0\ : std_logic;
signal \ADC_VDC.genclk.n21211_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21205\ : std_logic;
signal \ADC_VDC.genclk.t0on_13\ : std_logic;
signal \ADC_VDC.genclk.t0on_3\ : std_logic;
signal \ADC_VDC.genclk.t0on_5\ : std_logic;
signal \ADC_VDC.genclk.t0on_8\ : std_logic;
signal \ADC_VDC.genclk.n26_adj_1408\ : std_logic;
signal \ADC_VDC.genclk.t0on_14\ : std_logic;
signal \ADC_VDC.genclk.t0on_9\ : std_logic;
signal \ADC_VDC.genclk.t0on_15\ : std_logic;
signal \ADC_VDC.genclk.t0on_11\ : std_logic;
signal \ADC_VDC.genclk.n28_adj_1407\ : std_logic;
signal \ADC_VDC.genclk.t0on_12\ : std_logic;
signal \ADC_VDC.genclk.t0on_2\ : std_logic;
signal \ADC_VDC.genclk.t0on_7\ : std_logic;
signal \ADC_VDC.genclk.t0on_10\ : std_logic;
signal \ADC_VDC.genclk.n27_adj_1409\ : std_logic;
signal buf_data_vac_16 : std_logic;
signal buf_data_vac_20 : std_logic;
signal comm_buf_3_4 : std_logic;
signal buf_data_vac_23 : std_logic;
signal buf_data_vac_22 : std_logic;
signal buf_data_vac_21 : std_logic;
signal buf_data_vac_19 : std_logic;
signal buf_data_vac_18 : std_logic;
signal buf_data_vac_17 : std_logic;
signal n12152 : std_logic;
signal n14787 : std_logic;
signal \n1_cascade_\ : std_logic;
signal comm_buf_2_0 : std_logic;
signal comm_buf_3_0 : std_logic;
signal n2 : std_logic;
signal comm_buf_5_0 : std_logic;
signal n20970 : std_logic;
signal \n4_adj_1507_cascade_\ : std_logic;
signal n21980 : std_logic;
signal \n21116_cascade_\ : std_logic;
signal n10713 : std_logic;
signal n12_adj_1602 : std_logic;
signal buf_data_vac_8 : std_logic;
signal comm_buf_4_0 : std_logic;
signal buf_data_vac_15 : std_logic;
signal buf_data_vac_14 : std_logic;
signal buf_data_vac_13 : std_logic;
signal buf_data_vac_12 : std_logic;
signal comm_buf_4_4 : std_logic;
signal buf_data_vac_11 : std_logic;
signal buf_data_vac_10 : std_logic;
signal buf_data_vac_9 : std_logic;
signal n12194 : std_logic;
signal n14794 : std_logic;
signal \n1_adj_1589_cascade_\ : std_logic;
signal comm_buf_6_3 : std_logic;
signal \n21296_cascade_\ : std_logic;
signal n22154 : std_logic;
signal comm_buf_4_3 : std_logic;
signal comm_buf_5_3 : std_logic;
signal n4_adj_1591 : std_logic;
signal comm_buf_3_3 : std_logic;
signal comm_buf_2_3 : std_logic;
signal n2_adj_1590 : std_logic;
signal \n21102_cascade_\ : std_logic;
signal n21_adj_1618 : std_logic;
signal n16_adj_1599 : std_logic;
signal data_idxvec_6 : std_logic;
signal buf_data_iac_14 : std_logic;
signal \n26_adj_1505_cascade_\ : std_logic;
signal \n20930_cascade_\ : std_logic;
signal \n21962_cascade_\ : std_logic;
signal \n21965_cascade_\ : std_logic;
signal buf_adcdata_vdc_14 : std_logic;
signal buf_adcdata_vac_14 : std_logic;
signal \buf_readRTD_6\ : std_logic;
signal \n19_cascade_\ : std_logic;
signal n20954 : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal n20929 : std_logic;
signal comm_buf_1_3 : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal \n20884_cascade_\ : std_logic;
signal n20878 : std_logic;
signal \n22124_cascade_\ : std_logic;
signal n22127 : std_logic;
signal data_idxvec_3 : std_logic;
signal buf_data_iac_11 : std_logic;
signal \n26_adj_1514_cascade_\ : std_logic;
signal n20885 : std_logic;
signal \buf_readRTD_3\ : std_logic;
signal n20879 : std_logic;
signal buf_adcdata_vac_11 : std_logic;
signal buf_adcdata_vdc_11 : std_logic;
signal n19_adj_1513 : std_logic;
signal \n22178_cascade_\ : std_logic;
signal \n22181_cascade_\ : std_logic;
signal \n30_adj_1511_cascade_\ : std_logic;
signal data_idxvec_4 : std_logic;
signal n26_adj_1510 : std_logic;
signal n19_adj_1509 : std_logic;
signal \buf_readRTD_4\ : std_logic;
signal buf_adcdata_iac_12 : std_logic;
signal \n22010_cascade_\ : std_logic;
signal n16_adj_1508 : std_logic;
signal n22013 : std_logic;
signal \n12441_cascade_\ : std_logic;
signal \n8_adj_1567_cascade_\ : std_logic;
signal data_index_1 : std_logic;
signal n11835 : std_logic;
signal n16763 : std_logic;
signal buf_dds1_1 : std_logic;
signal buf_adcdata_iac_14 : std_logic;
signal n16 : std_logic;
signal n20953 : std_logic;
signal n10614 : std_logic;
signal n12312 : std_logic;
signal \VDC_RNG0\ : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal n12383 : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal n14 : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n18_adj_1611 : std_logic;
signal data_index_4 : std_logic;
signal n7_adj_1560 : std_logic;
signal n8_adj_1561 : std_logic;
signal \data_index_9_N_216_4\ : std_logic;
signal n8_adj_1565 : std_logic;
signal n7_adj_1564 : std_logic;
signal \data_index_9_N_216_2\ : std_logic;
signal n14_adj_1573 : std_logic;
signal n14_adj_1572 : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal n22_adj_1620 : std_logic;
signal n9_adj_1415 : std_logic;
signal n14_adj_1570 : std_logic;
signal n21048 : std_logic;
signal n10_adj_1613 : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal n19498 : std_logic;
signal n19499 : std_logic;
signal n19500 : std_logic;
signal n19501 : std_logic;
signal n19502 : std_logic;
signal n10 : std_logic;
signal n19503 : std_logic;
signal n19504 : std_logic;
signal \INVdds0_mclkcnt_i7_3783__i0C_net\ : std_logic;
signal secclk_cnt_0 : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal secclk_cnt_1 : std_logic;
signal n19509 : std_logic;
signal secclk_cnt_2 : std_logic;
signal n19510 : std_logic;
signal secclk_cnt_3 : std_logic;
signal n19511 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n19512 : std_logic;
signal secclk_cnt_5 : std_logic;
signal n19513 : std_logic;
signal secclk_cnt_6 : std_logic;
signal n19514 : std_logic;
signal secclk_cnt_7 : std_logic;
signal n19515 : std_logic;
signal n19516 : std_logic;
signal secclk_cnt_8 : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal secclk_cnt_9 : std_logic;
signal n19517 : std_logic;
signal secclk_cnt_10 : std_logic;
signal n19518 : std_logic;
signal secclk_cnt_11 : std_logic;
signal n19519 : std_logic;
signal secclk_cnt_12 : std_logic;
signal n19520 : std_logic;
signal secclk_cnt_13 : std_logic;
signal n19521 : std_logic;
signal secclk_cnt_14 : std_logic;
signal n19522 : std_logic;
signal secclk_cnt_15 : std_logic;
signal n19523 : std_logic;
signal n19524 : std_logic;
signal secclk_cnt_16 : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal secclk_cnt_17 : std_logic;
signal n19525 : std_logic;
signal secclk_cnt_18 : std_logic;
signal n19526 : std_logic;
signal secclk_cnt_19 : std_logic;
signal n19527 : std_logic;
signal secclk_cnt_20 : std_logic;
signal n19528 : std_logic;
signal secclk_cnt_21 : std_logic;
signal n19529 : std_logic;
signal n19530 : std_logic;
signal secclk_cnt_22 : std_logic;
signal n14731 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal \ADC_VDC.genclk.div_state_1\ : std_logic;
signal \VDC_CLK\ : std_logic;
signal \INVADC_VDC.genclk.t_clk_24C_net\ : std_logic;
signal \n21506_cascade_\ : std_logic;
signal n21067 : std_logic;
signal n23_adj_1538 : std_logic;
signal n22028 : std_logic;
signal buf_adcdata_iac_20 : std_logic;
signal buf_dds0_12 : std_logic;
signal \n22088_cascade_\ : std_logic;
signal buf_dds1_12 : std_logic;
signal \n22091_cascade_\ : std_logic;
signal n22205 : std_logic;
signal n22031 : std_logic;
signal \n20844_cascade_\ : std_logic;
signal comm_rx_buf_4 : std_logic;
signal \n30_adj_1539_cascade_\ : std_logic;
signal comm_cmd_7 : std_logic;
signal \n20621_cascade_\ : std_logic;
signal \n25_adj_1619_cascade_\ : std_logic;
signal \comm_spi.n16869\ : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal n7_adj_1609 : std_logic;
signal buf_dds1_11 : std_logic;
signal buf_dds0_11 : std_logic;
signal buf_adcdata_iac_19 : std_logic;
signal n22082 : std_logic;
signal data_idxvec_11 : std_logic;
signal buf_data_iac_19 : std_logic;
signal \n26_adj_1541_cascade_\ : std_logic;
signal \n20837_cascade_\ : std_logic;
signal n22085 : std_logic;
signal \n22094_cascade_\ : std_logic;
signal n20828 : std_logic;
signal comm_rx_buf_3 : std_logic;
signal \n22097_cascade_\ : std_logic;
signal flagcntwd : std_logic;
signal n11406 : std_logic;
signal \n12242_cascade_\ : std_logic;
signal \n20599_cascade_\ : std_logic;
signal n5 : std_logic;
signal \IAC_FLT1\ : std_logic;
signal eis_state_1 : std_logic;
signal buf_data_iac_8 : std_logic;
signal data_idxvec_12 : std_logic;
signal n20983 : std_logic;
signal n12397 : std_logic;
signal \VAC_OSR0\ : std_logic;
signal n21046 : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal n19_adj_1487 : std_logic;
signal \buf_readRTD_0\ : std_logic;
signal data_idxvec_0 : std_logic;
signal n20973 : std_logic;
signal \n26_cascade_\ : std_logic;
signal n21998 : std_logic;
signal n16_adj_1488 : std_logic;
signal n22004 : std_logic;
signal \n22007_cascade_\ : std_logic;
signal n22001 : std_logic;
signal \n30_adj_1486_cascade_\ : std_logic;
signal comm_buf_1_0 : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal eis_start : std_logic;
signal n21992 : std_logic;
signal data_idxvec_8 : std_logic;
signal buf_data_iac_16 : std_logic;
signal \n20917_cascade_\ : std_logic;
signal n21995 : std_logic;
signal \n20919_cascade_\ : std_logic;
signal n22043 : std_logic;
signal n22019 : std_logic;
signal \n22220_cascade_\ : std_logic;
signal \n22223_cascade_\ : std_logic;
signal comm_buf_0_0 : std_logic;
signal \iac_raw_buf_N_737\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal n19354 : std_logic;
signal n19355 : std_logic;
signal n19356 : std_logic;
signal n19357 : std_logic;
signal n19358 : std_logic;
signal n19359 : std_logic;
signal n19360 : std_logic;
signal n19361 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal n19362 : std_logic;
signal n19363 : std_logic;
signal n19364 : std_logic;
signal n19365 : std_logic;
signal n19366 : std_logic;
signal n19367 : std_logic;
signal n19368 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal n13473 : std_logic;
signal n14663 : std_logic;
signal data_cntvec_14 : std_logic;
signal data_cntvec_11 : std_logic;
signal req_data_cnt_14 : std_logic;
signal n8828 : std_logic;
signal \n8_adj_1559_cascade_\ : std_logic;
signal \data_index_9_N_216_6\ : std_logic;
signal n8_adj_1567 : std_logic;
signal n7_adj_1566 : std_logic;
signal \data_index_9_N_216_1\ : std_logic;
signal data_cntvec_12 : std_logic;
signal data_cntvec_10 : std_logic;
signal req_data_cnt_12 : std_logic;
signal req_data_cnt_10 : std_logic;
signal n8_adj_1559 : std_logic;
signal n7_adj_1558 : std_logic;
signal data_index_6 : std_logic;
signal \comm_spi.data_tx_7__N_771\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal n19505 : std_logic;
signal n19506 : std_logic;
signal n19507 : std_logic;
signal n19508 : std_logic;
signal clk_cnt_0 : std_logic;
signal clk_cnt_4 : std_logic;
signal clk_cnt_1 : std_logic;
signal clk_cnt_3 : std_logic;
signal \n6_cascade_\ : std_logic;
signal clk_cnt_2 : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal dds0_mclkcnt_3 : std_logic;
signal dds0_mclkcnt_5 : std_logic;
signal dds0_mclkcnt_1 : std_logic;
signal dds0_mclkcnt_4 : std_logic;
signal dds0_mclkcnt_2 : std_logic;
signal dds0_mclkcnt_0 : std_logic;
signal \n12_cascade_\ : std_logic;
signal dds0_mclkcnt_7 : std_logic;
signal n20543 : std_logic;
signal \n20543_cascade_\ : std_logic;
signal dds0_mclkcnt_6 : std_logic;
signal \INVdds0_mclk_304C_net\ : std_logic;
signal buf_data_iac_22 : std_logic;
signal n21038 : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal \INVcomm_spi.bit_cnt_3778__i3C_net\ : std_logic;
signal n30_adj_1529 : std_logic;
signal n22109 : std_logic;
signal n14766 : std_logic;
signal \n21199_cascade_\ : std_logic;
signal \n20681_cascade_\ : std_logic;
signal n20599 : std_logic;
signal \n12108_cascade_\ : std_logic;
signal n4_adj_1616 : std_logic;
signal n11977 : std_logic;
signal comm_buf_3_6 : std_logic;
signal comm_buf_2_6 : std_logic;
signal comm_buf_6_6 : std_logic;
signal \n21329_cascade_\ : std_logic;
signal \n21986_cascade_\ : std_logic;
signal n2_adj_1584 : std_logic;
signal comm_buf_0_6 : std_logic;
signal n1_adj_1583 : std_logic;
signal n20621 : std_logic;
signal \n7_cascade_\ : std_logic;
signal comm_buf_2_2 : std_logic;
signal comm_buf_3_2 : std_logic;
signal comm_buf_0_2 : std_logic;
signal \n22046_cascade_\ : std_logic;
signal comm_buf_5_2 : std_logic;
signal comm_buf_4_2 : std_logic;
signal comm_buf_6_2 : std_logic;
signal \n4_adj_1593_cascade_\ : std_logic;
signal n22049 : std_logic;
signal \n20801_cascade_\ : std_logic;
signal n20596 : std_logic;
signal n21094 : std_logic;
signal \n21092_cascade_\ : std_logic;
signal n20_adj_1610 : std_logic;
signal n20883 : std_logic;
signal \n20695_cascade_\ : std_logic;
signal n20881 : std_logic;
signal \n14545_cascade_\ : std_logic;
signal data_idxvec_1 : std_logic;
signal \n26_adj_1522_cascade_\ : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal \n22190_cascade_\ : std_logic;
signal \n22193_cascade_\ : std_logic;
signal \n30_adj_1523_cascade_\ : std_logic;
signal n19_adj_1520 : std_logic;
signal \buf_readRTD_1\ : std_logic;
signal \n22064_cascade_\ : std_logic;
signal n16_adj_1519 : std_logic;
signal n22067 : std_logic;
signal \buf_readRTD_5\ : std_logic;
signal buf_adcdata_iac_13 : std_logic;
signal \n22142_cascade_\ : std_logic;
signal n16_adj_1496 : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal n22145 : std_logic;
signal \n22133_cascade_\ : std_logic;
signal \n30_adj_1499_cascade_\ : std_logic;
signal data_idxvec_5 : std_logic;
signal \n26_adj_1498_cascade_\ : std_logic;
signal n22130 : std_logic;
signal data_cntvec_8 : std_logic;
signal data_cntvec_13 : std_logic;
signal \n19_adj_1597_cascade_\ : std_logic;
signal \n29_adj_1635_cascade_\ : std_logic;
signal n16_adj_1623 : std_logic;
signal req_data_cnt_8 : std_logic;
signal n10534 : std_logic;
signal n20798 : std_logic;
signal n22061 : std_logic;
signal n14730 : std_logic;
signal \clk_RTD\ : std_logic;
signal n23 : std_logic;
signal n21_adj_1521 : std_logic;
signal \n22_adj_1568_cascade_\ : std_logic;
signal n30_adj_1641 : std_logic;
signal data_idxvec_9 : std_logic;
signal buf_data_iac_17 : std_logic;
signal \n20812_cascade_\ : std_logic;
signal comm_buf_0_3 : std_logic;
signal \SELIRNG1\ : std_logic;
signal comm_buf_0_4 : std_logic;
signal n14_adj_1571 : std_logic;
signal n14_adj_1549 : std_logic;
signal n20814 : std_logic;
signal n22025 : std_logic;
signal \n22232_cascade_\ : std_logic;
signal n22235 : std_logic;
signal buf_adcdata_vdc_17 : std_logic;
signal buf_adcdata_vac_17 : std_logic;
signal n22226 : std_logic;
signal n22229 : std_logic;
signal \DDS_RNG_0\ : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal n22037 : std_logic;
signal buf_dds1_7 : std_logic;
signal buf_dds0_7 : std_logic;
signal req_data_cnt_11 : std_logic;
signal n23_adj_1540 : std_logic;
signal n20836 : std_logic;
signal n14_adj_1545 : std_logic;
signal n11931 : std_logic;
signal \n21073_cascade_\ : std_logic;
signal \n21072_cascade_\ : std_logic;
signal \clk_16MHz\ : std_logic;
signal dds0_mclk : std_logic;
signal buf_control_6 : std_logic;
signal \DDS_MCLK\ : std_logic;
signal buf_adcdata_iac_15 : std_logic;
signal n16_adj_1503 : std_logic;
signal n20797 : std_logic;
signal eis_stop : std_logic;
signal n22034 : std_logic;
signal \SIG_DDS.bit_cnt_1\ : std_logic;
signal \SIG_DDS.bit_cnt_2\ : std_logic;
signal \SIG_DDS.bit_cnt_3\ : std_logic;
signal trig_dds0 : std_logic;
signal n14900 : std_logic;
signal bit_cnt_0 : std_logic;
signal tmp_buf_15 : std_logic;
signal \DDS_MOSI\ : std_logic;
signal \DDS_CS\ : std_logic;
signal \SIG_DDS.n9_adj_1394\ : std_logic;
signal buf_data_iac_20 : std_logic;
signal n20984 : std_logic;
signal n17738 : std_logic;
signal n14146 : std_logic;
signal \comm_state_3_N_436_2\ : std_logic;
signal \n15_cascade_\ : std_logic;
signal n12_adj_1649 : std_logic;
signal comm_buf_4_1 : std_logic;
signal comm_buf_5_1 : std_logic;
signal \n4_adj_1595_cascade_\ : std_logic;
signal comm_buf_2_1 : std_logic;
signal comm_buf_3_1 : std_logic;
signal comm_buf_0_1 : std_logic;
signal \n22052_cascade_\ : std_logic;
signal comm_buf_1_1 : std_logic;
signal n20807 : std_logic;
signal \n22055_cascade_\ : std_logic;
signal comm_buf_5_5 : std_logic;
signal comm_buf_3_5 : std_logic;
signal \n17404_cascade_\ : std_logic;
signal \n20951_cascade_\ : std_logic;
signal comm_rx_buf_1 : std_logic;
signal comm_buf_6_1 : std_logic;
signal \n4_adj_1598_cascade_\ : std_logic;
signal n20573 : std_logic;
signal \comm_state_3_N_420_3\ : std_logic;
signal \n1272_cascade_\ : std_logic;
signal comm_buf_4_5 : std_logic;
signal n22175 : std_logic;
signal n20551 : std_logic;
signal n11420 : std_logic;
signal \n20551_cascade_\ : std_logic;
signal n20717 : std_logic;
signal n20575 : std_logic;
signal n20962 : std_logic;
signal n14545 : std_logic;
signal n22238 : std_logic;
signal \n2_adj_1575_cascade_\ : std_logic;
signal \n22241_cascade_\ : std_logic;
signal n8_adj_1576 : std_logic;
signal n1272 : std_logic;
signal n20697 : std_logic;
signal n4_adj_1614 : std_logic;
signal n20668 : std_logic;
signal n11866 : std_logic;
signal n14753 : std_logic;
signal n8_adj_1530 : std_logic;
signal comm_buf_3_7 : std_logic;
signal comm_buf_2_7 : std_logic;
signal \n2_adj_1581_cascade_\ : std_logic;
signal n11503 : std_logic;
signal n14815 : std_logic;
signal comm_buf_0_7 : std_logic;
signal n1_adj_1580 : std_logic;
signal comm_buf_5_7 : std_logic;
signal comm_buf_4_7 : std_logic;
signal n20966 : std_logic;
signal \n4_adj_1582_cascade_\ : std_logic;
signal n21968 : std_logic;
signal comm_buf_1_5 : std_logic;
signal buf_data_iac_9 : std_logic;
signal n21270 : std_logic;
signal n9 : std_logic;
signal n20663 : std_logic;
signal \n12467_cascade_\ : std_logic;
signal n14_adj_1533 : std_logic;
signal data_cntvec_6 : std_logic;
signal data_cntvec_0 : std_logic;
signal req_data_cnt_0 : std_logic;
signal n17 : std_logic;
signal n16_adj_1515 : std_logic;
signal comm_buf_0_5 : std_logic;
signal req_data_cnt_6 : std_logic;
signal req_data_cnt_2 : std_logic;
signal \n22208_cascade_\ : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal n21959 : std_logic;
signal \n22211_cascade_\ : std_logic;
signal comm_rx_buf_2 : std_logic;
signal \n30_adj_1518_cascade_\ : std_logic;
signal comm_buf_1_2 : std_logic;
signal n12047 : std_logic;
signal n14773 : std_logic;
signal n19_adj_1516 : std_logic;
signal \buf_readRTD_2\ : std_logic;
signal n21956 : std_logic;
signal data_idxvec_2 : std_logic;
signal data_cntvec_2 : std_logic;
signal n26_adj_1517 : std_logic;
signal n14_adj_1550 : std_logic;
signal n14_adj_1544 : std_logic;
signal data_cntvec_1 : std_logic;
signal data_cntvec_4 : std_logic;
signal req_data_cnt_4 : std_logic;
signal req_data_cnt_1 : std_logic;
signal n18 : std_logic;
signal buf_adcdata_vdc_13 : std_logic;
signal buf_adcdata_vac_13 : std_logic;
signal n19_adj_1497 : std_logic;
signal n14_adj_1579 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal n23_adj_1527 : std_logic;
signal data_cntvec_5 : std_logic;
signal data_cntvec_3 : std_logic;
signal req_data_cnt_3 : std_logic;
signal n20_adj_1596 : std_logic;
signal comm_buf_1_7 : std_logic;
signal n14_adj_1546 : std_logic;
signal \n14_adj_1546_cascade_\ : std_logic;
signal n14_adj_1577 : std_logic;
signal req_data_cnt_13 : std_logic;
signal data_cntvec_9 : std_logic;
signal req_data_cnt_15 : std_logic;
signal data_cntvec_15 : std_logic;
signal n24 : std_logic;
signal n14_adj_1574 : std_logic;
signal req_data_cnt_9 : std_logic;
signal n12467 : std_logic;
signal n14_adj_1578 : std_logic;
signal req_data_cnt_5 : std_logic;
signal n9321 : std_logic;
signal n12441 : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal data_idxvec_7 : std_logic;
signal data_cntvec_7 : std_logic;
signal buf_data_iac_15 : std_logic;
signal \n26_adj_1500_cascade_\ : std_logic;
signal \n20810_cascade_\ : std_logic;
signal n22058 : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal req_data_cnt_7 : std_logic;
signal n20809 : std_logic;
signal comm_cmd_2 : std_logic;
signal comm_cmd_3 : std_logic;
signal comm_cmd_1 : std_logic;
signal comm_length_1 : std_logic;
signal comm_length_2 : std_logic;
signal comm_length_0 : std_logic;
signal n4 : std_logic;
signal n14671 : std_logic;
signal \SIG_DDS.n21331\ : std_logic;
signal \SIG_DDS.n10\ : std_logic;
signal \SIG_DDS.n9\ : std_logic;
signal dds_state_0 : std_logic;
signal dds_state_2 : std_logic;
signal dds_state_1 : std_logic;
signal \DDS_SCK\ : std_logic;
signal wdtick_flag : std_logic;
signal buf_control_0 : std_logic;
signal \CONT_SD\ : std_logic;
signal n20608 : std_logic;
signal n23_adj_1501 : std_logic;
signal \n21_adj_1600_cascade_\ : std_logic;
signal n17485 : std_logic;
signal n18_adj_1633 : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.n22667\ : std_logic;
signal \comm_spi.n14630\ : std_logic;
signal \comm_spi.n22667_cascade_\ : std_logic;
signal comm_rx_buf_0 : std_logic;
signal \comm_rx_buf_0_cascade_\ : std_logic;
signal comm_buf_6_0 : std_logic;
signal comm_index_2 : std_logic;
signal comm_buf_2_5 : std_logic;
signal comm_index_1 : std_logic;
signal n22172 : std_logic;
signal comm_rx_buf_5 : std_logic;
signal comm_buf_6_5 : std_logic;
signal \n2369_cascade_\ : std_logic;
signal \n21130_cascade_\ : std_logic;
signal n14_adj_1506 : std_logic;
signal n3 : std_logic;
signal n20681 : std_logic;
signal \n3_cascade_\ : std_logic;
signal n2369 : std_logic;
signal n19655 : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal comm_data_vld : std_logic;
signal n21129 : std_logic;
signal n20740 : std_logic;
signal \n11363_cascade_\ : std_logic;
signal n12242 : std_logic;
signal n12235 : std_logic;
signal n11869 : std_logic;
signal n11876 : std_logic;
signal comm_rx_buf_7 : std_logic;
signal n12244 : std_logic;
signal comm_buf_6_7 : std_logic;
signal \THERMOSTAT\ : std_logic;
signal buf_control_7 : std_logic;
signal n11935 : std_logic;
signal n19904 : std_logic;
signal comm_buf_1_4 : std_logic;
signal n14_adj_1548 : std_logic;
signal cmd_rdadctmp_20_adj_1430 : std_logic;
signal comm_buf_1_6 : std_logic;
signal comm_state_2 : std_logic;
signal n14_adj_1547 : std_logic;
signal buf_adcdata_iac_8 : std_logic;
signal cmd_rdadctmp_16_adj_1434 : std_logic;
signal n12663 : std_logic;
signal cmd_rdadctmp_18_adj_1432 : std_logic;
signal buf_adcdata_iac_10 : std_logic;
signal cmd_rdadctmp_19_adj_1431 : std_logic;
signal buf_adcdata_iac_11 : std_logic;
signal n20584 : std_logic;
signal adc_state_0_adj_1418 : std_logic;
signal cmd_rdadctmp_17_adj_1433 : std_logic;
signal buf_adcdata_iac_9 : std_logic;
signal buf_data_iac_12 : std_logic;
signal n21230 : std_logic;
signal buf_data_iac_13 : std_logic;
signal n21297 : std_logic;
signal \comm_spi.DOUT_7__N_747\ : std_logic;
signal comm_state_3 : std_logic;
signal n11377 : std_logic;
signal \comm_spi.data_tx_7__N_770\ : std_logic;
signal comm_buf_5_6 : std_logic;
signal comm_buf_4_6 : std_logic;
signal comm_index_0 : std_logic;
signal n4_adj_1585 : std_logic;
signal comm_state_1 : std_logic;
signal comm_state_0 : std_logic;
signal n9270 : std_logic;
signal \comm_spi.n22670\ : std_logic;
signal \comm_spi.n14631\ : std_logic;
signal \comm_spi.n14616\ : std_logic;
signal \comm_spi.n14617\ : std_logic;
signal \INVcomm_spi.imiso_83_12208_12209_setC_net\ : std_logic;
signal comm_tx_buf_2 : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.DOUT_7__N_748\ : std_logic;
signal \comm_spi.imosi_N_753\ : std_logic;
signal \comm_spi.data_tx_7__N_790\ : std_logic;
signal \comm_spi.n22685\ : std_logic;
signal \comm_spi.data_tx_7__N_772\ : std_logic;
signal \comm_spi.n14634\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal \comm_spi.data_tx_7__N_773\ : std_logic;
signal \comm_spi.n22682\ : std_logic;
signal \comm_spi.n14638\ : std_logic;
signal \comm_spi.n14639\ : std_logic;
signal \comm_spi.data_tx_7__N_787\ : std_logic;
signal comm_tx_buf_3 : std_logic;
signal comm_tx_buf_4 : std_logic;
signal comm_tx_buf_5 : std_logic;
signal \comm_spi.n22679\ : std_logic;
signal \comm_spi.n14642\ : std_logic;
signal \comm_spi.n14643\ : std_logic;
signal \comm_spi.data_tx_7__N_784\ : std_logic;
signal \comm_spi.data_tx_7__N_781\ : std_logic;
signal buf_data_iac_23 : std_logic;
signal n21204 : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \comm_spi.n14621\ : std_logic;
signal \INVcomm_spi.MISO_48_12202_12203_resetC_net\ : std_logic;
signal \comm_spi.n14626\ : std_logic;
signal \comm_spi.n14620\ : std_logic;
signal \INVcomm_spi.MISO_48_12202_12203_setC_net\ : std_logic;
signal comm_tx_buf_6 : std_logic;
signal \comm_spi.n14619\ : std_logic;
signal \comm_spi.n14627\ : std_logic;
signal \INVcomm_spi.imiso_83_12208_12209_resetC_net\ : std_logic;
signal \comm_spi.n14624\ : std_logic;
signal \comm_spi.n22661\ : std_logic;
signal \comm_spi.n14623\ : std_logic;
signal \comm_spi.data_tx_7__N_767\ : std_logic;
signal comm_tx_buf_7 : std_logic;
signal \comm_spi.data_tx_7__N_775\ : std_logic;
signal \comm_spi.n14635\ : std_logic;
signal \comm_spi.data_tx_7__N_793\ : std_logic;
signal \comm_spi.n22664\ : std_logic;
signal \comm_spi.n14612\ : std_logic;
signal \comm_spi.iclk_N_763\ : std_logic;
signal \comm_spi.n22688\ : std_logic;
signal comm_cmd_0 : std_logic;
signal buf_data_iac_10 : std_logic;
signal n21320 : std_logic;
signal \comm_spi.n14655\ : std_logic;
signal \comm_spi.data_tx_7__N_778\ : std_logic;
signal \comm_spi.n22673\ : std_logic;
signal \comm_spi.n14651\ : std_logic;
signal \comm_spi.n14654\ : std_logic;
signal \comm_spi.data_tx_7__N_768\ : std_logic;
signal \comm_spi.n22676\ : std_logic;
signal \comm_spi.n14646\ : std_logic;
signal \comm_spi.n14647\ : std_logic;
signal \comm_spi.n14650\ : std_logic;
signal \comm_spi.data_tx_7__N_769\ : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_754\ : std_logic;
signal \comm_spi.n14608\ : std_logic;
signal \comm_spi.data_tx_7__N_774\ : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.n14613\ : std_logic;
signal \clk_32MHz\ : std_logic;
signal \comm_spi.iclk_N_764\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \comm_spi.n14609\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal comm_clear : std_logic;
signal comm_tx_buf_0 : std_logic;
signal \comm_spi.data_tx_7__N_796\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VAC_DRDY_wire\ : std_logic;
signal \IAC_FLT1_wire\ : std_logic;
signal \DDS_SCK_wire\ : std_logic;
signal \ICE_IOR_166_wire\ : std_logic;
signal \ICE_IOR_119_wire\ : std_logic;
signal \DDS_MOSI_wire\ : std_logic;
signal \VAC_MISO_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \ICE_IOR_146_wire\ : std_logic;
signal \VDC_CLK_wire\ : std_logic;
signal \ICE_IOT_222_wire\ : std_logic;
signal \IAC_CS_wire\ : std_logic;
signal \ICE_IOL_18B_wire\ : std_logic;
signal \ICE_IOL_13A_wire\ : std_logic;
signal \ICE_IOB_81_wire\ : std_logic;
signal \VAC_OSR1_wire\ : std_logic;
signal \IAC_MOSI_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \ICE_IOL_4B_wire\ : std_logic;
signal \ICE_IOB_94_wire\ : std_logic;
signal \VAC_CS_wire\ : std_logic;
signal \VAC_CLK_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \ICE_IOR_167_wire\ : std_logic;
signal \ICE_IOR_118_wire\ : std_logic;
signal \RTD_SDO_wire\ : std_logic;
signal \IAC_OSR0_wire\ : std_logic;
signal \VDC_SCLK_wire\ : std_logic;
signal \VAC_FLT1_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_IOR_165_wire\ : std_logic;
signal \ICE_IOR_147_wire\ : std_logic;
signal \ICE_IOL_14A_wire\ : std_logic;
signal \ICE_IOL_13B_wire\ : std_logic;
signal \ICE_IOB_91_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_RNG_0_wire\ : std_logic;
signal \VDC_RNG0_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \ICE_IOR_152_wire\ : std_logic;
signal \ICE_IOL_12A_wire\ : std_logic;
signal \RTD_DRDY_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_IOT_177_wire\ : std_logic;
signal \ICE_IOR_141_wire\ : std_logic;
signal \ICE_IOB_102_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \IAC_MISO_wire\ : std_logic;
signal \VAC_OSR0_wire\ : std_logic;
signal \VAC_MOSI_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \ICE_IOR_148_wire\ : std_logic;
signal \STAT_COMM_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \ICE_IOR_161_wire\ : std_logic;
signal \ICE_IOB_95_wire\ : std_logic;
signal \ICE_IOB_82_wire\ : std_logic;
signal \ICE_IOB_104_wire\ : std_logic;
signal \IAC_CLK_wire\ : std_logic;
signal \DDS_CS_wire\ : std_logic;
signal \SELIRNG0_wire\ : std_logic;
signal \RTD_SDI_wire\ : std_logic;
signal \ICE_IOT_221_wire\ : std_logic;
signal \ICE_IOT_197_wire\ : std_logic;
signal \DDS_MCLK_wire\ : std_logic;
signal \RTD_SCLK_wire\ : std_logic;
signal \RTD_CS_wire\ : std_logic;
signal \ICE_IOR_137_wire\ : std_logic;
signal \IAC_OSR1_wire\ : std_logic;
signal \VAC_FLT0_wire\ : std_logic;
signal \ICE_IOR_144_wire\ : std_logic;
signal \ICE_IOR_128_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \IAC_SCLK_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \ICE_IOR_139_wire\ : std_logic;
signal \ICE_IOL_4A_wire\ : std_logic;
signal \VAC_SCLK_wire\ : std_logic;
signal \THERMOSTAT_wire\ : std_logic;
signal \ICE_IOR_164_wire\ : std_logic;
signal \ICE_IOB_103_wire\ : std_logic;
signal \OUT_SYNCCLK_wire\ : std_logic;
signal \AMPV_POW_wire\ : std_logic;
signal \VDC_SDO_wire\ : std_logic;
signal \ICE_IOT_174_wire\ : std_logic;
signal \ICE_IOR_140_wire\ : std_logic;
signal \ICE_IOB_96_wire\ : std_logic;
signal \CONT_SD_wire\ : std_logic;
signal \AC_ADC_SYNC_wire\ : std_logic;
signal \SELIRNG1_wire\ : std_logic;
signal \ICE_IOL_12B_wire\ : std_logic;
signal \ICE_IOR_160_wire\ : std_logic;
signal \ICE_IOR_136_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_IOT_198_wire\ : std_logic;
signal \ICE_IOT_173_wire\ : std_logic;
signal \IAC_DRDY_wire\ : std_logic;
signal \ICE_IOT_178_wire\ : std_logic;
signal \ICE_IOR_138_wire\ : std_logic;
signal \ICE_IOR_120_wire\ : std_logic;
signal \IAC_FLT0_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \VAC_DRDY_wire\ <= VAC_DRDY;
    IAC_FLT1 <= \IAC_FLT1_wire\;
    DDS_SCK <= \DDS_SCK_wire\;
    \ICE_IOR_166_wire\ <= ICE_IOR_166;
    \ICE_IOR_119_wire\ <= ICE_IOR_119;
    DDS_MOSI <= \DDS_MOSI_wire\;
    \VAC_MISO_wire\ <= VAC_MISO;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    \ICE_IOR_146_wire\ <= ICE_IOR_146;
    VDC_CLK <= \VDC_CLK_wire\;
    \ICE_IOT_222_wire\ <= ICE_IOT_222;
    IAC_CS <= \IAC_CS_wire\;
    \ICE_IOL_18B_wire\ <= ICE_IOL_18B;
    \ICE_IOL_13A_wire\ <= ICE_IOL_13A;
    \ICE_IOB_81_wire\ <= ICE_IOB_81;
    VAC_OSR1 <= \VAC_OSR1_wire\;
    IAC_MOSI <= \IAC_MOSI_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    \ICE_IOL_4B_wire\ <= ICE_IOL_4B;
    \ICE_IOB_94_wire\ <= ICE_IOB_94;
    VAC_CS <= \VAC_CS_wire\;
    VAC_CLK <= \VAC_CLK_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    \ICE_IOR_167_wire\ <= ICE_IOR_167;
    \ICE_IOR_118_wire\ <= ICE_IOR_118;
    \RTD_SDO_wire\ <= RTD_SDO;
    IAC_OSR0 <= \IAC_OSR0_wire\;
    VDC_SCLK <= \VDC_SCLK_wire\;
    VAC_FLT1 <= \VAC_FLT1_wire\;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_IOR_165_wire\ <= ICE_IOR_165;
    \ICE_IOR_147_wire\ <= ICE_IOR_147;
    \ICE_IOL_14A_wire\ <= ICE_IOL_14A;
    \ICE_IOL_13B_wire\ <= ICE_IOL_13B;
    \ICE_IOB_91_wire\ <= ICE_IOB_91;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_RNG_0 <= \DDS_RNG_0_wire\;
    VDC_RNG0 <= \VDC_RNG0_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    \ICE_IOR_152_wire\ <= ICE_IOR_152;
    \ICE_IOL_12A_wire\ <= ICE_IOL_12A;
    \RTD_DRDY_wire\ <= RTD_DRDY;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_IOT_177_wire\ <= ICE_IOT_177;
    \ICE_IOR_141_wire\ <= ICE_IOR_141;
    \ICE_IOB_102_wire\ <= ICE_IOB_102;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    \IAC_MISO_wire\ <= IAC_MISO;
    VAC_OSR0 <= \VAC_OSR0_wire\;
    VAC_MOSI <= \VAC_MOSI_wire\;
    TEST_LED <= \TEST_LED_wire\;
    \ICE_IOR_148_wire\ <= ICE_IOR_148;
    STAT_COMM <= \STAT_COMM_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    \ICE_IOR_161_wire\ <= ICE_IOR_161;
    \ICE_IOB_95_wire\ <= ICE_IOB_95;
    \ICE_IOB_82_wire\ <= ICE_IOB_82;
    \ICE_IOB_104_wire\ <= ICE_IOB_104;
    IAC_CLK <= \IAC_CLK_wire\;
    DDS_CS <= \DDS_CS_wire\;
    SELIRNG0 <= \SELIRNG0_wire\;
    RTD_SDI <= \RTD_SDI_wire\;
    \ICE_IOT_221_wire\ <= ICE_IOT_221;
    \ICE_IOT_197_wire\ <= ICE_IOT_197;
    DDS_MCLK <= \DDS_MCLK_wire\;
    RTD_SCLK <= \RTD_SCLK_wire\;
    RTD_CS <= \RTD_CS_wire\;
    \ICE_IOR_137_wire\ <= ICE_IOR_137;
    IAC_OSR1 <= \IAC_OSR1_wire\;
    VAC_FLT0 <= \VAC_FLT0_wire\;
    \ICE_IOR_144_wire\ <= ICE_IOR_144;
    \ICE_IOR_128_wire\ <= ICE_IOR_128;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    IAC_SCLK <= \IAC_SCLK_wire\;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    \ICE_IOR_139_wire\ <= ICE_IOR_139;
    \ICE_IOL_4A_wire\ <= ICE_IOL_4A;
    VAC_SCLK <= \VAC_SCLK_wire\;
    \THERMOSTAT_wire\ <= THERMOSTAT;
    \ICE_IOR_164_wire\ <= ICE_IOR_164;
    \ICE_IOB_103_wire\ <= ICE_IOB_103;
    OUT_SYNCCLK <= \OUT_SYNCCLK_wire\;
    AMPV_POW <= \AMPV_POW_wire\;
    \VDC_SDO_wire\ <= VDC_SDO;
    \ICE_IOT_174_wire\ <= ICE_IOT_174;
    \ICE_IOR_140_wire\ <= ICE_IOR_140;
    \ICE_IOB_96_wire\ <= ICE_IOB_96;
    CONT_SD <= \CONT_SD_wire\;
    AC_ADC_SYNC <= \AC_ADC_SYNC_wire\;
    SELIRNG1 <= \SELIRNG1_wire\;
    \ICE_IOL_12B_wire\ <= ICE_IOL_12B;
    \ICE_IOR_160_wire\ <= ICE_IOR_160;
    \ICE_IOR_136_wire\ <= ICE_IOR_136;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_IOT_198_wire\ <= ICE_IOT_198;
    \ICE_IOT_173_wire\ <= ICE_IOT_173;
    \IAC_DRDY_wire\ <= IAC_DRDY;
    \ICE_IOT_178_wire\ <= ICE_IOT_178;
    \ICE_IOR_138_wire\ <= ICE_IOR_138;
    \ICE_IOR_120_wire\ <= ICE_IOR_120;
    IAC_FLT0 <= \IAC_FLT0_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data_iac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(13);
    buf_data_vac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(9);
    buf_data_iac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(5);
    buf_data_vac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ <= '0'&\N__28217\&\N__25697\&\N__27800\&\N__42278\&\N__31142\&\N__38690\&\N__35978\&\N__39389\&\N__42152\&\N__27350\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ <= '0'&\N__30668\&\N__30776\&\N__29600\&\N__29708\&\N__29810\&\N__29924\&\N__30029\&\N__30143\&\N__30251\&\N__30359\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ <= '0'&'0'&\N__40913\&'0'&'0'&'0'&\N__29429\&'0'&'0'&'0'&\N__27455\&'0'&'0'&'0'&\N__29033\&'0';
    buf_data_iac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(13);
    buf_data_vac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(9);
    buf_data_iac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(5);
    buf_data_vac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ <= '0'&\N__28171\&\N__25660\&\N__27760\&\N__42238\&\N__31108\&\N__38653\&\N__35938\&\N__39352\&\N__42115\&\N__27313\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ <= '0'&\N__30631\&\N__30733\&\N__29563\&\N__29668\&\N__29776\&\N__29890\&\N__29998\&\N__30112\&\N__30214\&\N__30322\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ <= '0'&'0'&\N__52613\&'0'&'0'&'0'&\N__30833\&'0'&'0'&'0'&\N__52153\&'0'&'0'&'0'&\N__30524\&'0';
    buf_data_iac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(13);
    buf_data_vac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(9);
    buf_data_iac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(5);
    buf_data_vac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ <= '0'&\N__28235\&\N__25715\&\N__27818\&\N__42296\&\N__31160\&\N__38708\&\N__35996\&\N__39407\&\N__42170\&\N__27368\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ <= '0'&\N__30686\&\N__30794\&\N__29618\&\N__29726\&\N__29828\&\N__29942\&\N__30047\&\N__30161\&\N__30269\&\N__30377\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ <= '0'&'0'&\N__22892\&'0'&'0'&'0'&\N__25487\&'0'&'0'&'0'&\N__40382\&'0'&'0'&'0'&\N__21953\&'0';
    buf_data_iac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(13);
    buf_data_vac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(9);
    buf_data_iac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(5);
    buf_data_vac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ <= '0'&\N__28183\&\N__25672\&\N__27772\&\N__42250\&\N__31118\&\N__38665\&\N__35950\&\N__39364\&\N__42127\&\N__27325\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ <= '0'&\N__30643\&\N__30745\&\N__29575\&\N__29680\&\N__29786\&\N__29900\&\N__30005\&\N__30119\&\N__30226\&\N__30334\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ <= '0'&'0'&\N__53237\&'0'&'0'&'0'&\N__38294\&'0'&'0'&'0'&\N__51875\&'0'&'0'&'0'&\N__30473\&'0';
    buf_data_iac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(13);
    buf_data_vac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(9);
    buf_data_iac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(5);
    buf_data_vac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ <= '0'&\N__28241\&\N__25721\&\N__27824\&\N__42302\&\N__31166\&\N__38714\&\N__36002\&\N__39413\&\N__42176\&\N__27374\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ <= '0'&\N__30692\&\N__30800\&\N__29624\&\N__29732\&\N__29834\&\N__29948\&\N__30053\&\N__30167\&\N__30275\&\N__30383\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ <= '0'&'0'&\N__22859\&'0'&'0'&'0'&\N__22277\&'0'&'0'&'0'&\N__36820\&'0'&'0'&'0'&\N__31967\&'0';
    buf_data_iac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(13);
    buf_data_vac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(9);
    buf_data_iac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(5);
    buf_data_vac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ <= '0'&\N__28195\&\N__25679\&\N__27782\&\N__42260\&\N__31124\&\N__38672\&\N__35960\&\N__39371\&\N__42134\&\N__27332\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ <= '0'&\N__30650\&\N__30757\&\N__29582\&\N__29690\&\N__29792\&\N__29906\&\N__30011\&\N__30125\&\N__30233\&\N__30341\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ <= '0'&'0'&\N__43579\&'0'&'0'&'0'&\N__46649\&'0'&'0'&'0'&\N__38165\&'0'&'0'&'0'&\N__35603\&'0';
    buf_data_iac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(13);
    buf_data_vac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(9);
    buf_data_iac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(5);
    buf_data_vac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ <= '0'&\N__28192\&\N__25663\&\N__27769\&\N__42247\&\N__31105\&\N__38656\&\N__35947\&\N__39355\&\N__42118\&\N__27316\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ <= '0'&\N__30634\&\N__30748\&\N__29566\&\N__29677\&\N__29773\&\N__29887\&\N__29989\&\N__30103\&\N__30217\&\N__30325\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ <= '0'&'0'&\N__25865\&'0'&'0'&'0'&\N__21977\&'0'&'0'&'0'&\N__21869\&'0'&'0'&'0'&\N__21893\&'0';
    buf_data_iac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(13);
    buf_data_vac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(9);
    buf_data_iac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(5);
    buf_data_vac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ <= '0'&\N__28205\&\N__25685\&\N__27788\&\N__42266\&\N__31130\&\N__38678\&\N__35966\&\N__39377\&\N__42140\&\N__27338\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ <= '0'&\N__30656\&\N__30764\&\N__29588\&\N__29696\&\N__29798\&\N__29912\&\N__30017\&\N__30131\&\N__30239\&\N__30347\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ <= '0'&'0'&\N__44959\&'0'&'0'&'0'&\N__29324\&'0'&'0'&'0'&\N__38366\&'0'&'0'&'0'&\N__38084\&'0';
    buf_data_iac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(13);
    buf_data_vac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(9);
    buf_data_iac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(5);
    buf_data_vac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ <= '0'&\N__28204\&\N__25675\&\N__27781\&\N__42259\&\N__31117\&\N__38668\&\N__35959\&\N__39367\&\N__42130\&\N__27328\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ <= '0'&\N__30646\&\N__30760\&\N__29578\&\N__29689\&\N__29785\&\N__29899\&\N__30001\&\N__30115\&\N__30229\&\N__30337\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ <= '0'&'0'&\N__23630\&'0'&'0'&'0'&\N__23654\&'0'&'0'&'0'&\N__23771\&'0'&'0'&'0'&\N__23591\&'0';
    buf_data_iac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(13);
    buf_data_vac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(9);
    buf_data_iac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(5);
    buf_data_vac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ <= '0'&\N__28229\&\N__25709\&\N__27812\&\N__42290\&\N__31154\&\N__38702\&\N__35990\&\N__39401\&\N__42164\&\N__27362\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ <= '0'&\N__30680\&\N__30788\&\N__29612\&\N__29720\&\N__29822\&\N__29936\&\N__30041\&\N__30155\&\N__30263\&\N__30371\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ <= '0'&'0'&\N__28472\&'0'&'0'&'0'&\N__28802\&'0'&'0'&'0'&\N__28592\&'0'&'0'&'0'&\N__28619\&'0';
    buf_data_iac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(13);
    buf_data_vac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(9);
    buf_data_iac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(5);
    buf_data_vac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ <= '0'&\N__28211\&\N__25691\&\N__27794\&\N__42272\&\N__31136\&\N__38684\&\N__35972\&\N__39383\&\N__42146\&\N__27344\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ <= '0'&\N__30662\&\N__30770\&\N__29594\&\N__29702\&\N__29804\&\N__29918\&\N__30023\&\N__30137\&\N__30245\&\N__30353\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ <= '0'&'0'&\N__25556\&'0'&'0'&'0'&\N__43967\&'0'&'0'&'0'&\N__22793\&'0'&'0'&'0'&\N__30410\&'0';
    buf_data_iac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(13);
    buf_data_vac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(9);
    buf_data_iac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(5);
    buf_data_vac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ <= '0'&\N__28223\&\N__25703\&\N__27806\&\N__42284\&\N__31148\&\N__38696\&\N__35984\&\N__39395\&\N__42158\&\N__27356\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ <= '0'&\N__30674\&\N__30782\&\N__29606\&\N__29714\&\N__29816\&\N__29930\&\N__30035\&\N__30149\&\N__30257\&\N__30365\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ <= '0'&'0'&\N__28913\&'0'&'0'&'0'&\N__34745\&'0'&'0'&'0'&\N__34070\&'0'&'0'&'0'&\N__33964\&'0';

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__19205\,
            RESETB => \N__57232\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \clk_16MHz\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \iac_raw_buf_vac_raw_buf_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57931\,
            RE => \N__57187\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            WE => \N__35539\
        );

    \iac_raw_buf_vac_raw_buf_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57982\,
            RE => \N__57379\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            WE => \N__35568\
        );

    \iac_raw_buf_vac_raw_buf_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57858\,
            RE => \N__57147\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            WE => \N__35567\
        );

    \iac_raw_buf_vac_raw_buf_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57980\,
            RE => \N__57320\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            WE => \N__35566\
        );

    \iac_raw_buf_vac_raw_buf_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57837\,
            RE => \N__57167\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            WE => \N__35570\
        );

    \iac_raw_buf_vac_raw_buf_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57977\,
            RE => \N__57319\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            WE => \N__35554\
        );

    \iac_raw_buf_vac_raw_buf_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57848\,
            RE => \N__57380\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            WE => \N__35558\
        );

    \iac_raw_buf_vac_raw_buf_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57968\,
            RE => \N__57238\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            WE => \N__35546\
        );

    \iac_raw_buf_vac_raw_buf_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57827\,
            RE => \N__57318\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            WE => \N__35569\
        );

    \iac_raw_buf_vac_raw_buf_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57877\,
            RE => \N__57148\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            WE => \N__35562\
        );

    \iac_raw_buf_vac_raw_buf_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57954\,
            RE => \N__57236\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            WE => \N__35506\
        );

    \iac_raw_buf_vac_raw_buf_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__57905\,
            RE => \N__57185\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            WE => \N__35550\
        );

    \ipInertedIOPad_VAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59184\,
            DIN => \N__59183\,
            DOUT => \N__59182\,
            PACKAGEPIN => \VAC_DRDY_wire\
        );

    \ipInertedIOPad_VAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59184\,
            PADOUT => \N__59183\,
            PADIN => \N__59182\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59175\,
            DIN => \N__59174\,
            DOUT => \N__59173\,
            PACKAGEPIN => \IAC_FLT1_wire\
        );

    \ipInertedIOPad_IAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59175\,
            PADOUT => \N__59174\,
            PADIN => \N__59173\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41093\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59166\,
            DIN => \N__59165\,
            DOUT => \N__59164\,
            PACKAGEPIN => \DDS_SCK_wire\
        );

    \ipInertedIOPad_DDS_SCK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59166\,
            PADOUT => \N__59165\,
            PADIN => \N__59164\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__50039\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_166_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59157\,
            DIN => \N__59156\,
            DOUT => \N__59155\,
            PACKAGEPIN => \ICE_IOR_166_wire\
        );

    \ipInertedIOPad_ICE_IOR_166_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59157\,
            PADOUT => \N__59156\,
            PADIN => \N__59155\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_119_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59148\,
            DIN => \N__59147\,
            DOUT => \N__59146\,
            PACKAGEPIN => \ICE_IOR_119_wire\
        );

    \ipInertedIOPad_ICE_IOR_119_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59148\,
            PADOUT => \N__59147\,
            PADIN => \N__59146\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59139\,
            DIN => \N__59138\,
            DOUT => \N__59137\,
            PACKAGEPIN => \DDS_MOSI_wire\
        );

    \ipInertedIOPad_DDS_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59139\,
            PADOUT => \N__59138\,
            PADIN => \N__59137\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44705\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59130\,
            DIN => \N__59129\,
            DOUT => \N__59128\,
            PACKAGEPIN => \VAC_MISO_wire\
        );

    \ipInertedIOPad_VAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59130\,
            PADOUT => \N__59129\,
            PADIN => \N__59128\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59121\,
            DIN => \N__59120\,
            DOUT => \N__59119\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59121\,
            PADOUT => \N__59120\,
            PADIN => \N__59119\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21722\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_146_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59112\,
            DIN => \N__59111\,
            DOUT => \N__59110\,
            PACKAGEPIN => \ICE_IOR_146_wire\
        );

    \ipInertedIOPad_ICE_IOR_146_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59112\,
            PADOUT => \N__59111\,
            PADIN => \N__59110\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59103\,
            DIN => \N__59102\,
            DOUT => \N__59101\,
            PACKAGEPIN => \VDC_CLK_wire\
        );

    \ipInertedIOPad_VDC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59103\,
            PADOUT => \N__59102\,
            PADIN => \N__59101\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__40089\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_222_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59094\,
            DIN => \N__59093\,
            DOUT => \N__59092\,
            PACKAGEPIN => \ICE_IOT_222_wire\
        );

    \ipInertedIOPad_ICE_IOT_222_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59094\,
            PADOUT => \N__59093\,
            PADIN => \N__59092\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59085\,
            DIN => \N__59084\,
            DOUT => \N__59083\,
            PACKAGEPIN => \IAC_CS_wire\
        );

    \ipInertedIOPad_IAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59085\,
            PADOUT => \N__59084\,
            PADIN => \N__59083\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20621\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_18B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59076\,
            DIN => \N__59075\,
            DOUT => \N__59074\,
            PACKAGEPIN => \ICE_IOL_18B_wire\
        );

    \ipInertedIOPad_ICE_IOL_18B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59076\,
            PADOUT => \N__59075\,
            PADIN => \N__59074\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59067\,
            DIN => \N__59066\,
            DOUT => \N__59065\,
            PACKAGEPIN => \ICE_IOL_13A_wire\
        );

    \ipInertedIOPad_ICE_IOL_13A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59067\,
            PADOUT => \N__59066\,
            PADIN => \N__59065\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_81_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59058\,
            DIN => \N__59057\,
            DOUT => \N__59056\,
            PACKAGEPIN => \ICE_IOB_81_wire\
        );

    \ipInertedIOPad_ICE_IOB_81_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59058\,
            PADOUT => \N__59057\,
            PADIN => \N__59056\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59049\,
            DIN => \N__59048\,
            DOUT => \N__59047\,
            PACKAGEPIN => \VAC_OSR1_wire\
        );

    \ipInertedIOPad_VAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59049\,
            PADOUT => \N__59048\,
            PADIN => \N__59047\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22913\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59040\,
            DIN => \N__59039\,
            DOUT => \N__59038\,
            PACKAGEPIN => \IAC_MOSI_wire\
        );

    \ipInertedIOPad_IAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59040\,
            PADOUT => \N__59039\,
            PADIN => \N__59038\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59031\,
            DIN => \N__59030\,
            DOUT => \N__59029\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59031\,
            PADOUT => \N__59030\,
            PADIN => \N__59029\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19841\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59022\,
            DIN => \N__59021\,
            DOUT => \N__59020\,
            PACKAGEPIN => \ICE_IOL_4B_wire\
        );

    \ipInertedIOPad_ICE_IOL_4B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59022\,
            PADOUT => \N__59021\,
            PADIN => \N__59020\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_94_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59013\,
            DIN => \N__59012\,
            DOUT => \N__59011\,
            PACKAGEPIN => \ICE_IOB_94_wire\
        );

    \ipInertedIOPad_ICE_IOB_94_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59013\,
            PADOUT => \N__59012\,
            PADIN => \N__59011\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59004\,
            DIN => \N__59003\,
            DOUT => \N__59002\,
            PACKAGEPIN => \VAC_CS_wire\
        );

    \ipInertedIOPad_VAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59004\,
            PADOUT => \N__59003\,
            PADIN => \N__59002\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19448\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58995\,
            DIN => \N__58994\,
            DOUT => \N__58993\,
            PACKAGEPIN => \VAC_CLK_wire\
        );

    \ipInertedIOPad_VAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58995\,
            PADOUT => \N__58994\,
            PADIN => \N__58993\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23068\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58986\,
            DIN => \N__58985\,
            DOUT => \N__58984\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58986\,
            PADOUT => \N__58985\,
            PADIN => \N__58984\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_167_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58977\,
            DIN => \N__58976\,
            DOUT => \N__58975\,
            PACKAGEPIN => \ICE_IOR_167_wire\
        );

    \ipInertedIOPad_ICE_IOR_167_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58977\,
            PADOUT => \N__58976\,
            PADIN => \N__58975\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_118_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58968\,
            DIN => \N__58967\,
            DOUT => \N__58966\,
            PACKAGEPIN => \ICE_IOR_118_wire\
        );

    \ipInertedIOPad_ICE_IOR_118_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58968\,
            PADOUT => \N__58967\,
            PADIN => \N__58966\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDO_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58959\,
            DIN => \N__58958\,
            DOUT => \N__58957\,
            PACKAGEPIN => \RTD_SDO_wire\
        );

    \ipInertedIOPad_RTD_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58959\,
            PADOUT => \N__58958\,
            PADIN => \N__58957\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58950\,
            DIN => \N__58949\,
            DOUT => \N__58948\,
            PACKAGEPIN => \IAC_OSR0_wire\
        );

    \ipInertedIOPad_IAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58950\,
            PADOUT => \N__58949\,
            PADIN => \N__58948\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22760\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58941\,
            DIN => \N__58940\,
            DOUT => \N__58939\,
            PACKAGEPIN => \VDC_SCLK_wire\
        );

    \ipInertedIOPad_VDC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58941\,
            PADOUT => \N__58940\,
            PADIN => \N__58939\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21092\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58932\,
            DIN => \N__58931\,
            DOUT => \N__58930\,
            PACKAGEPIN => \VAC_FLT1_wire\
        );

    \ipInertedIOPad_VAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58932\,
            PADOUT => \N__58931\,
            PADIN => \N__58930\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22835\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58923\,
            DIN => \N__58922\,
            DOUT => \N__58921\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58923\,
            PADOUT => \N__58922\,
            PADIN => \N__58921\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_165_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58914\,
            DIN => \N__58913\,
            DOUT => \N__58912\,
            PACKAGEPIN => \ICE_IOR_165_wire\
        );

    \ipInertedIOPad_ICE_IOR_165_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58914\,
            PADOUT => \N__58913\,
            PADIN => \N__58912\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_147_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58905\,
            DIN => \N__58904\,
            DOUT => \N__58903\,
            PACKAGEPIN => \ICE_IOR_147_wire\
        );

    \ipInertedIOPad_ICE_IOR_147_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58905\,
            PADOUT => \N__58904\,
            PADIN => \N__58903\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_14A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58896\,
            DIN => \N__58895\,
            DOUT => \N__58894\,
            PACKAGEPIN => \ICE_IOL_14A_wire\
        );

    \ipInertedIOPad_ICE_IOL_14A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58896\,
            PADOUT => \N__58895\,
            PADIN => \N__58894\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58887\,
            DIN => \N__58886\,
            DOUT => \N__58885\,
            PACKAGEPIN => \ICE_IOL_13B_wire\
        );

    \ipInertedIOPad_ICE_IOL_13B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58887\,
            PADOUT => \N__58886\,
            PADIN => \N__58885\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_91_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58878\,
            DIN => \N__58877\,
            DOUT => \N__58876\,
            PACKAGEPIN => \ICE_IOB_91_wire\
        );

    \ipInertedIOPad_ICE_IOB_91_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58878\,
            PADOUT => \N__58877\,
            PADIN => \N__58876\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58869\,
            DIN => \N__58868\,
            DOUT => \N__58867\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58869\,
            PADOUT => \N__58868\,
            PADIN => \N__58867\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_RNG_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58860\,
            DIN => \N__58859\,
            DOUT => \N__58858\,
            PACKAGEPIN => \DDS_RNG_0_wire\
        );

    \ipInertedIOPad_DDS_RNG_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58860\,
            PADOUT => \N__58859\,
            PADIN => \N__58858\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44660\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_RNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58851\,
            DIN => \N__58850\,
            DOUT => \N__58849\,
            PACKAGEPIN => \VDC_RNG0_wire\
        );

    \ipInertedIOPad_VDC_RNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58851\,
            PADOUT => \N__58850\,
            PADIN => \N__58849\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39035\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58842\,
            DIN => \N__58841\,
            DOUT => \N__58840\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58842\,
            PADOUT => \N__58841\,
            PADIN => \N__58840\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_152_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58833\,
            DIN => \N__58832\,
            DOUT => \N__58831\,
            PACKAGEPIN => \ICE_IOR_152_wire\
        );

    \ipInertedIOPad_ICE_IOR_152_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58833\,
            PADOUT => \N__58832\,
            PADIN => \N__58831\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58824\,
            DIN => \N__58823\,
            DOUT => \N__58822\,
            PACKAGEPIN => \ICE_IOL_12A_wire\
        );

    \ipInertedIOPad_ICE_IOL_12A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58824\,
            PADOUT => \N__58823\,
            PADIN => \N__58822\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_DRDY_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58815\,
            DIN => \N__58814\,
            DOUT => \N__58813\,
            PACKAGEPIN => \RTD_DRDY_wire\
        );

    \ipInertedIOPad_RTD_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58815\,
            PADOUT => \N__58814\,
            PADIN => \N__58813\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58806\,
            DIN => \N__58805\,
            DOUT => \N__58804\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58806\,
            PADOUT => \N__58805\,
            PADIN => \N__58804\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__55565\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_177_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58797\,
            DIN => \N__58796\,
            DOUT => \N__58795\,
            PACKAGEPIN => \ICE_IOT_177_wire\
        );

    \ipInertedIOPad_ICE_IOT_177_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58797\,
            PADOUT => \N__58796\,
            PADIN => \N__58795\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_141_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58788\,
            DIN => \N__58787\,
            DOUT => \N__58786\,
            PACKAGEPIN => \ICE_IOR_141_wire\
        );

    \ipInertedIOPad_ICE_IOR_141_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58788\,
            PADOUT => \N__58787\,
            PADIN => \N__58786\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_102_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58779\,
            DIN => \N__58778\,
            DOUT => \N__58777\,
            PACKAGEPIN => \ICE_IOB_102_wire\
        );

    \ipInertedIOPad_ICE_IOB_102_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58779\,
            PADOUT => \N__58778\,
            PADIN => \N__58777\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58770\,
            DIN => \N__58769\,
            DOUT => \N__58768\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58770\,
            PADOUT => \N__58769\,
            PADIN => \N__58768\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58761\,
            DIN => \N__58760\,
            DOUT => \N__58759\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58761\,
            PADOUT => \N__58760\,
            PADIN => \N__58759\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27971\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58752\,
            DIN => \N__58751\,
            DOUT => \N__58750\,
            PACKAGEPIN => \IAC_MISO_wire\
        );

    \ipInertedIOPad_IAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58752\,
            PADOUT => \N__58751\,
            PADIN => \N__58750\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58743\,
            DIN => \N__58742\,
            DOUT => \N__58741\,
            PACKAGEPIN => \VAC_OSR0_wire\
        );

    \ipInertedIOPad_VAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58743\,
            PADOUT => \N__58742\,
            PADIN => \N__58741\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41339\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58734\,
            DIN => \N__58733\,
            DOUT => \N__58732\,
            PACKAGEPIN => \VAC_MOSI_wire\
        );

    \ipInertedIOPad_VAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58734\,
            PADOUT => \N__58733\,
            PADIN => \N__58732\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58725\,
            DIN => \N__58724\,
            DOUT => \N__58723\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58725\,
            PADOUT => \N__58724\,
            PADIN => \N__58723\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32741\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_148_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58716\,
            DIN => \N__58715\,
            DOUT => \N__58714\,
            PACKAGEPIN => \ICE_IOR_148_wire\
        );

    \ipInertedIOPad_ICE_IOR_148_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58716\,
            PADOUT => \N__58715\,
            PADIN => \N__58714\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_STAT_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58707\,
            DIN => \N__58706\,
            DOUT => \N__58705\,
            PACKAGEPIN => \STAT_COMM_wire\
        );

    \ipInertedIOPad_STAT_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58707\,
            PADOUT => \N__58706\,
            PADIN => \N__58705\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19190\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58698\,
            DIN => \N__58697\,
            DOUT => \N__58696\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58698\,
            PADOUT => \N__58697\,
            PADIN => \N__58696\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_161_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58689\,
            DIN => \N__58688\,
            DOUT => \N__58687\,
            PACKAGEPIN => \ICE_IOR_161_wire\
        );

    \ipInertedIOPad_ICE_IOR_161_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58689\,
            PADOUT => \N__58688\,
            PADIN => \N__58687\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_95_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58680\,
            DIN => \N__58679\,
            DOUT => \N__58678\,
            PACKAGEPIN => \ICE_IOB_95_wire\
        );

    \ipInertedIOPad_ICE_IOB_95_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58680\,
            PADOUT => \N__58679\,
            PADIN => \N__58678\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_82_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58671\,
            DIN => \N__58670\,
            DOUT => \N__58669\,
            PACKAGEPIN => \ICE_IOB_82_wire\
        );

    \ipInertedIOPad_ICE_IOB_82_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58671\,
            PADOUT => \N__58670\,
            PADIN => \N__58669\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_104_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58662\,
            DIN => \N__58661\,
            DOUT => \N__58660\,
            PACKAGEPIN => \ICE_IOB_104_wire\
        );

    \ipInertedIOPad_ICE_IOB_104_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58662\,
            PADOUT => \N__58661\,
            PADIN => \N__58660\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58653\,
            DIN => \N__58652\,
            DOUT => \N__58651\,
            PACKAGEPIN => \IAC_CLK_wire\
        );

    \ipInertedIOPad_IAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58653\,
            PADOUT => \N__58652\,
            PADIN => \N__58651\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23075\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58644\,
            DIN => \N__58643\,
            DOUT => \N__58642\,
            PACKAGEPIN => \DDS_CS_wire\
        );

    \ipInertedIOPad_DDS_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58644\,
            PADOUT => \N__58643\,
            PADIN => \N__58642\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__45278\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58635\,
            DIN => \N__58634\,
            DOUT => \N__58633\,
            PACKAGEPIN => \SELIRNG0_wire\
        );

    \ipInertedIOPad_SELIRNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58635\,
            PADOUT => \N__58634\,
            PADIN => \N__58633\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23024\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58626\,
            DIN => \N__58625\,
            DOUT => \N__58624\,
            PACKAGEPIN => \RTD_SDI_wire\
        );

    \ipInertedIOPad_RTD_SDI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58626\,
            PADOUT => \N__58625\,
            PADIN => \N__58624\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20348\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_221_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58617\,
            DIN => \N__58616\,
            DOUT => \N__58615\,
            PACKAGEPIN => \ICE_IOT_221_wire\
        );

    \ipInertedIOPad_ICE_IOT_221_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58617\,
            PADOUT => \N__58616\,
            PADIN => \N__58615\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_197_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58608\,
            DIN => \N__58607\,
            DOUT => \N__58606\,
            PACKAGEPIN => \ICE_IOT_197_wire\
        );

    \ipInertedIOPad_ICE_IOT_197_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58608\,
            PADOUT => \N__58607\,
            PADIN => \N__58606\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58599\,
            DIN => \N__58598\,
            DOUT => \N__58597\,
            PACKAGEPIN => \DDS_MCLK_wire\
        );

    \ipInertedIOPad_DDS_MCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58599\,
            PADOUT => \N__58598\,
            PADIN => \N__58597\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44984\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58590\,
            DIN => \N__58589\,
            DOUT => \N__58588\,
            PACKAGEPIN => \RTD_SCLK_wire\
        );

    \ipInertedIOPad_RTD_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58590\,
            PADOUT => \N__58589\,
            PADIN => \N__58588\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22205\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58581\,
            DIN => \N__58580\,
            DOUT => \N__58579\,
            PACKAGEPIN => \RTD_CS_wire\
        );

    \ipInertedIOPad_RTD_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58581\,
            PADOUT => \N__58580\,
            PADIN => \N__58579\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22355\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_137_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58572\,
            DIN => \N__58571\,
            DOUT => \N__58570\,
            PACKAGEPIN => \ICE_IOR_137_wire\
        );

    \ipInertedIOPad_ICE_IOR_137_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58572\,
            PADOUT => \N__58571\,
            PADIN => \N__58570\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58563\,
            DIN => \N__58562\,
            DOUT => \N__58561\,
            PACKAGEPIN => \IAC_OSR1_wire\
        );

    \ipInertedIOPad_IAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58563\,
            PADOUT => \N__58562\,
            PADIN => \N__58561\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27713\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58554\,
            DIN => \N__58553\,
            DOUT => \N__58552\,
            PACKAGEPIN => \VAC_FLT0_wire\
        );

    \ipInertedIOPad_VAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58554\,
            PADOUT => \N__58553\,
            PADIN => \N__58552\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36869\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_144_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58545\,
            DIN => \N__58544\,
            DOUT => \N__58543\,
            PACKAGEPIN => \ICE_IOR_144_wire\
        );

    \ipInertedIOPad_ICE_IOR_144_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58545\,
            PADOUT => \N__58544\,
            PADIN => \N__58543\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_128_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58536\,
            DIN => \N__58535\,
            DOUT => \N__58534\,
            PACKAGEPIN => \ICE_IOR_128_wire\
        );

    \ipInertedIOPad_ICE_IOR_128_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58536\,
            PADOUT => \N__58535\,
            PADIN => \N__58534\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58527\,
            DIN => \N__58526\,
            DOUT => \N__58525\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58527\,
            PADOUT => \N__58526\,
            PADIN => \N__58525\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_1\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58518\,
            DIN => \N__58517\,
            DOUT => \N__58516\,
            PACKAGEPIN => \IAC_SCLK_wire\
        );

    \ipInertedIOPad_IAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58518\,
            PADOUT => \N__58517\,
            PADIN => \N__58516\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20021\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58509\,
            DIN => \N__58508\,
            DOUT => \N__58507\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58509\,
            PADOUT => \N__58508\,
            PADIN => \N__58507\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \EIS_SYNCCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_139_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58500\,
            DIN => \N__58499\,
            DOUT => \N__58498\,
            PACKAGEPIN => \ICE_IOR_139_wire\
        );

    \ipInertedIOPad_ICE_IOR_139_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58500\,
            PADOUT => \N__58499\,
            PADIN => \N__58498\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58491\,
            DIN => \N__58490\,
            DOUT => \N__58489\,
            PACKAGEPIN => \ICE_IOL_4A_wire\
        );

    \ipInertedIOPad_ICE_IOL_4A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58491\,
            PADOUT => \N__58490\,
            PADIN => \N__58489\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58482\,
            DIN => \N__58481\,
            DOUT => \N__58480\,
            PACKAGEPIN => \VAC_SCLK_wire\
        );

    \ipInertedIOPad_VAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58482\,
            PADOUT => \N__58481\,
            PADIN => \N__58480\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19478\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_THERMOSTAT_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58473\,
            DIN => \N__58472\,
            DOUT => \N__58471\,
            PACKAGEPIN => \THERMOSTAT_wire\
        );

    \ipInertedIOPad_THERMOSTAT_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58473\,
            PADOUT => \N__58472\,
            PADIN => \N__58471\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \THERMOSTAT\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_164_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58464\,
            DIN => \N__58463\,
            DOUT => \N__58462\,
            PACKAGEPIN => \ICE_IOR_164_wire\
        );

    \ipInertedIOPad_ICE_IOR_164_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58464\,
            PADOUT => \N__58463\,
            PADIN => \N__58462\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_103_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58455\,
            DIN => \N__58454\,
            DOUT => \N__58453\,
            PACKAGEPIN => \ICE_IOB_103_wire\
        );

    \ipInertedIOPad_ICE_IOB_103_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58455\,
            PADOUT => \N__58454\,
            PADIN => \N__58453\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_OUT_SYNCCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58446\,
            DIN => \N__58445\,
            DOUT => \N__58444\,
            PACKAGEPIN => \OUT_SYNCCLK_wire\
        );

    \ipInertedIOPad_OUT_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58446\,
            PADOUT => \N__58445\,
            PADIN => \N__58444\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31346\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AMPV_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58437\,
            DIN => \N__58436\,
            DOUT => \N__58435\,
            PACKAGEPIN => \AMPV_POW_wire\
        );

    \ipInertedIOPad_AMPV_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58437\,
            PADOUT => \N__58436\,
            PADIN => \N__58435\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30956\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SDO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58428\,
            DIN => \N__58427\,
            DOUT => \N__58426\,
            PACKAGEPIN => \VDC_SDO_wire\
        );

    \ipInertedIOPad_VDC_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58428\,
            PADOUT => \N__58427\,
            PADIN => \N__58426\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VDC_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_174_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58419\,
            DIN => \N__58418\,
            DOUT => \N__58417\,
            PACKAGEPIN => \ICE_IOT_174_wire\
        );

    \ipInertedIOPad_ICE_IOT_174_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58419\,
            PADOUT => \N__58418\,
            PADIN => \N__58417\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_140_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58410\,
            DIN => \N__58409\,
            DOUT => \N__58408\,
            PACKAGEPIN => \ICE_IOR_140_wire\
        );

    \ipInertedIOPad_ICE_IOR_140_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58410\,
            PADOUT => \N__58409\,
            PADIN => \N__58408\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_96_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58401\,
            DIN => \N__58400\,
            DOUT => \N__58399\,
            PACKAGEPIN => \ICE_IOB_96_wire\
        );

    \ipInertedIOPad_ICE_IOB_96_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58401\,
            PADOUT => \N__58400\,
            PADIN => \N__58399\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CONT_SD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58392\,
            DIN => \N__58391\,
            DOUT => \N__58390\,
            PACKAGEPIN => \CONT_SD_wire\
        );

    \ipInertedIOPad_CONT_SD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58392\,
            PADOUT => \N__58391\,
            PADIN => \N__58390\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__49952\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AC_ADC_SYNC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58383\,
            DIN => \N__58382\,
            DOUT => \N__58381\,
            PACKAGEPIN => \AC_ADC_SYNC_wire\
        );

    \ipInertedIOPad_AC_ADC_SYNC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58383\,
            PADOUT => \N__58382\,
            PADIN => \N__58381\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25766\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58374\,
            DIN => \N__58373\,
            DOUT => \N__58372\,
            PACKAGEPIN => \SELIRNG1_wire\
        );

    \ipInertedIOPad_SELIRNG1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58374\,
            PADOUT => \N__58373\,
            PADIN => \N__58372\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44201\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58365\,
            DIN => \N__58364\,
            DOUT => \N__58363\,
            PACKAGEPIN => \ICE_IOL_12B_wire\
        );

    \ipInertedIOPad_ICE_IOL_12B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58365\,
            PADOUT => \N__58364\,
            PADIN => \N__58363\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_160_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58356\,
            DIN => \N__58355\,
            DOUT => \N__58354\,
            PACKAGEPIN => \ICE_IOR_160_wire\
        );

    \ipInertedIOPad_ICE_IOR_160_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58356\,
            PADOUT => \N__58355\,
            PADIN => \N__58354\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_136_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58347\,
            DIN => \N__58346\,
            DOUT => \N__58345\,
            PACKAGEPIN => \ICE_IOR_136_wire\
        );

    \ipInertedIOPad_ICE_IOR_136_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58347\,
            PADOUT => \N__58346\,
            PADIN => \N__58345\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58338\,
            DIN => \N__58337\,
            DOUT => \N__58336\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58338\,
            PADOUT => \N__58337\,
            PADIN => \N__58336\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20738\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_198_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58329\,
            DIN => \N__58328\,
            DOUT => \N__58327\,
            PACKAGEPIN => \ICE_IOT_198_wire\
        );

    \ipInertedIOPad_ICE_IOT_198_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58329\,
            PADOUT => \N__58328\,
            PADIN => \N__58327\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_173_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58320\,
            DIN => \N__58319\,
            DOUT => \N__58318\,
            PACKAGEPIN => \ICE_IOT_173_wire\
        );

    \ipInertedIOPad_ICE_IOT_173_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58320\,
            PADOUT => \N__58319\,
            PADIN => \N__58318\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58311\,
            DIN => \N__58310\,
            DOUT => \N__58309\,
            PACKAGEPIN => \IAC_DRDY_wire\
        );

    \ipInertedIOPad_IAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58311\,
            PADOUT => \N__58310\,
            PADIN => \N__58309\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_178_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58302\,
            DIN => \N__58301\,
            DOUT => \N__58300\,
            PACKAGEPIN => \ICE_IOT_178_wire\
        );

    \ipInertedIOPad_ICE_IOT_178_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58302\,
            PADOUT => \N__58301\,
            PADIN => \N__58300\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_138_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58293\,
            DIN => \N__58292\,
            DOUT => \N__58291\,
            PACKAGEPIN => \ICE_IOR_138_wire\
        );

    \ipInertedIOPad_ICE_IOR_138_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58293\,
            PADOUT => \N__58292\,
            PADIN => \N__58291\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_120_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58284\,
            DIN => \N__58283\,
            DOUT => \N__58282\,
            PACKAGEPIN => \ICE_IOR_120_wire\
        );

    \ipInertedIOPad_ICE_IOR_120_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58284\,
            PADOUT => \N__58283\,
            PADIN => \N__58282\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58275\,
            DIN => \N__58274\,
            DOUT => \N__58273\,
            PACKAGEPIN => \IAC_FLT0_wire\
        );

    \ipInertedIOPad_IAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58275\,
            PADOUT => \N__58274\,
            PADIN => \N__58273\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27416\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58266\,
            DIN => \N__58265\,
            DOUT => \N__58264\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58266\,
            PADOUT => \N__58265\,
            PADIN => \N__58264\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19883\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__14593\ : SRMux
    port map (
            O => \N__58247\,
            I => \N__58244\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__58244\,
            I => \comm_spi.data_tx_7__N_768\
        );

    \I__14591\ : InMux
    port map (
            O => \N__58241\,
            I => \N__58238\
        );

    \I__14590\ : LocalMux
    port map (
            O => \N__58238\,
            I => \N__58234\
        );

    \I__14589\ : InMux
    port map (
            O => \N__58237\,
            I => \N__58231\
        );

    \I__14588\ : Span4Mux_v
    port map (
            O => \N__58234\,
            I => \N__58228\
        );

    \I__14587\ : LocalMux
    port map (
            O => \N__58231\,
            I => \N__58225\
        );

    \I__14586\ : Span4Mux_v
    port map (
            O => \N__58228\,
            I => \N__58221\
        );

    \I__14585\ : Span4Mux_v
    port map (
            O => \N__58225\,
            I => \N__58218\
        );

    \I__14584\ : InMux
    port map (
            O => \N__58224\,
            I => \N__58215\
        );

    \I__14583\ : Odrv4
    port map (
            O => \N__58221\,
            I => \comm_spi.n22676\
        );

    \I__14582\ : Odrv4
    port map (
            O => \N__58218\,
            I => \comm_spi.n22676\
        );

    \I__14581\ : LocalMux
    port map (
            O => \N__58215\,
            I => \comm_spi.n22676\
        );

    \I__14580\ : InMux
    port map (
            O => \N__58208\,
            I => \N__58204\
        );

    \I__14579\ : InMux
    port map (
            O => \N__58207\,
            I => \N__58201\
        );

    \I__14578\ : LocalMux
    port map (
            O => \N__58204\,
            I => \N__58198\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__58201\,
            I => \comm_spi.n14646\
        );

    \I__14576\ : Odrv4
    port map (
            O => \N__58198\,
            I => \comm_spi.n14646\
        );

    \I__14575\ : InMux
    port map (
            O => \N__58193\,
            I => \N__58189\
        );

    \I__14574\ : InMux
    port map (
            O => \N__58192\,
            I => \N__58186\
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__58189\,
            I => \comm_spi.n14647\
        );

    \I__14572\ : LocalMux
    port map (
            O => \N__58186\,
            I => \comm_spi.n14647\
        );

    \I__14571\ : InMux
    port map (
            O => \N__58181\,
            I => \N__58178\
        );

    \I__14570\ : LocalMux
    port map (
            O => \N__58178\,
            I => \N__58174\
        );

    \I__14569\ : InMux
    port map (
            O => \N__58177\,
            I => \N__58171\
        );

    \I__14568\ : Odrv4
    port map (
            O => \N__58174\,
            I => \comm_spi.n14650\
        );

    \I__14567\ : LocalMux
    port map (
            O => \N__58171\,
            I => \comm_spi.n14650\
        );

    \I__14566\ : SRMux
    port map (
            O => \N__58166\,
            I => \N__58163\
        );

    \I__14565\ : LocalMux
    port map (
            O => \N__58163\,
            I => \N__58160\
        );

    \I__14564\ : Span4Mux_h
    port map (
            O => \N__58160\,
            I => \N__58157\
        );

    \I__14563\ : Odrv4
    port map (
            O => \N__58157\,
            I => \comm_spi.data_tx_7__N_769\
        );

    \I__14562\ : InMux
    port map (
            O => \N__58154\,
            I => \N__58149\
        );

    \I__14561\ : InMux
    port map (
            O => \N__58153\,
            I => \N__58146\
        );

    \I__14560\ : InMux
    port map (
            O => \N__58152\,
            I => \N__58143\
        );

    \I__14559\ : LocalMux
    port map (
            O => \N__58149\,
            I => \N__58136\
        );

    \I__14558\ : LocalMux
    port map (
            O => \N__58146\,
            I => \N__58136\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__58143\,
            I => \N__58136\
        );

    \I__14556\ : Span4Mux_v
    port map (
            O => \N__58136\,
            I => \N__58132\
        );

    \I__14555\ : InMux
    port map (
            O => \N__58135\,
            I => \N__58129\
        );

    \I__14554\ : Span4Mux_h
    port map (
            O => \N__58132\,
            I => \N__58125\
        );

    \I__14553\ : LocalMux
    port map (
            O => \N__58129\,
            I => \N__58122\
        );

    \I__14552\ : InMux
    port map (
            O => \N__58128\,
            I => \N__58119\
        );

    \I__14551\ : Sp12to4
    port map (
            O => \N__58125\,
            I => \N__58116\
        );

    \I__14550\ : Span4Mux_h
    port map (
            O => \N__58122\,
            I => \N__58113\
        );

    \I__14549\ : LocalMux
    port map (
            O => \N__58119\,
            I => \N__58110\
        );

    \I__14548\ : Span12Mux_s6_h
    port map (
            O => \N__58116\,
            I => \N__58103\
        );

    \I__14547\ : Sp12to4
    port map (
            O => \N__58113\,
            I => \N__58103\
        );

    \I__14546\ : Span12Mux_v
    port map (
            O => \N__58110\,
            I => \N__58103\
        );

    \I__14545\ : Span12Mux_v
    port map (
            O => \N__58103\,
            I => \N__58100\
        );

    \I__14544\ : Odrv12
    port map (
            O => \N__58100\,
            I => \ICE_SPI_MOSI\
        );

    \I__14543\ : SRMux
    port map (
            O => \N__58097\,
            I => \N__58094\
        );

    \I__14542\ : LocalMux
    port map (
            O => \N__58094\,
            I => \N__58091\
        );

    \I__14541\ : Span4Mux_h
    port map (
            O => \N__58091\,
            I => \N__58088\
        );

    \I__14540\ : Odrv4
    port map (
            O => \N__58088\,
            I => \comm_spi.imosi_N_754\
        );

    \I__14539\ : InMux
    port map (
            O => \N__58085\,
            I => \N__58081\
        );

    \I__14538\ : InMux
    port map (
            O => \N__58084\,
            I => \N__58078\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__58081\,
            I => \N__58073\
        );

    \I__14536\ : LocalMux
    port map (
            O => \N__58078\,
            I => \N__58073\
        );

    \I__14535\ : Span4Mux_h
    port map (
            O => \N__58073\,
            I => \N__58070\
        );

    \I__14534\ : Odrv4
    port map (
            O => \N__58070\,
            I => \comm_spi.n14608\
        );

    \I__14533\ : SRMux
    port map (
            O => \N__58067\,
            I => \N__58064\
        );

    \I__14532\ : LocalMux
    port map (
            O => \N__58064\,
            I => \N__58061\
        );

    \I__14531\ : Span4Mux_h
    port map (
            O => \N__58061\,
            I => \N__58058\
        );

    \I__14530\ : Odrv4
    port map (
            O => \N__58058\,
            I => \comm_spi.data_tx_7__N_774\
        );

    \I__14529\ : InMux
    port map (
            O => \N__58055\,
            I => \N__58051\
        );

    \I__14528\ : InMux
    port map (
            O => \N__58054\,
            I => \N__58048\
        );

    \I__14527\ : LocalMux
    port map (
            O => \N__58051\,
            I => \N__58045\
        );

    \I__14526\ : LocalMux
    port map (
            O => \N__58048\,
            I => \N__58042\
        );

    \I__14525\ : Span4Mux_v
    port map (
            O => \N__58045\,
            I => \N__58038\
        );

    \I__14524\ : Span4Mux_v
    port map (
            O => \N__58042\,
            I => \N__58035\
        );

    \I__14523\ : InMux
    port map (
            O => \N__58041\,
            I => \N__58032\
        );

    \I__14522\ : Span4Mux_h
    port map (
            O => \N__58038\,
            I => \N__58025\
        );

    \I__14521\ : Span4Mux_v
    port map (
            O => \N__58035\,
            I => \N__58025\
        );

    \I__14520\ : LocalMux
    port map (
            O => \N__58032\,
            I => \N__58022\
        );

    \I__14519\ : InMux
    port map (
            O => \N__58031\,
            I => \N__58019\
        );

    \I__14518\ : InMux
    port map (
            O => \N__58030\,
            I => \N__58016\
        );

    \I__14517\ : Sp12to4
    port map (
            O => \N__58025\,
            I => \N__58013\
        );

    \I__14516\ : Sp12to4
    port map (
            O => \N__58022\,
            I => \N__58006\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__58019\,
            I => \N__58006\
        );

    \I__14514\ : LocalMux
    port map (
            O => \N__58016\,
            I => \N__58006\
        );

    \I__14513\ : Span12Mux_s8_h
    port map (
            O => \N__58013\,
            I => \N__58001\
        );

    \I__14512\ : Span12Mux_v
    port map (
            O => \N__58006\,
            I => \N__58001\
        );

    \I__14511\ : Span12Mux_v
    port map (
            O => \N__58001\,
            I => \N__57998\
        );

    \I__14510\ : Odrv12
    port map (
            O => \N__57998\,
            I => \ICE_SPI_SCLK\
        );

    \I__14509\ : InMux
    port map (
            O => \N__57995\,
            I => \N__57992\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__57992\,
            I => \N__57989\
        );

    \I__14507\ : Span4Mux_v
    port map (
            O => \N__57989\,
            I => \N__57986\
        );

    \I__14506\ : Odrv4
    port map (
            O => \N__57986\,
            I => \comm_spi.n14613\
        );

    \I__14505\ : ClkMux
    port map (
            O => \N__57983\,
            I => \N__57443\
        );

    \I__14504\ : ClkMux
    port map (
            O => \N__57982\,
            I => \N__57443\
        );

    \I__14503\ : ClkMux
    port map (
            O => \N__57981\,
            I => \N__57443\
        );

    \I__14502\ : ClkMux
    port map (
            O => \N__57980\,
            I => \N__57443\
        );

    \I__14501\ : ClkMux
    port map (
            O => \N__57979\,
            I => \N__57443\
        );

    \I__14500\ : ClkMux
    port map (
            O => \N__57978\,
            I => \N__57443\
        );

    \I__14499\ : ClkMux
    port map (
            O => \N__57977\,
            I => \N__57443\
        );

    \I__14498\ : ClkMux
    port map (
            O => \N__57976\,
            I => \N__57443\
        );

    \I__14497\ : ClkMux
    port map (
            O => \N__57975\,
            I => \N__57443\
        );

    \I__14496\ : ClkMux
    port map (
            O => \N__57974\,
            I => \N__57443\
        );

    \I__14495\ : ClkMux
    port map (
            O => \N__57973\,
            I => \N__57443\
        );

    \I__14494\ : ClkMux
    port map (
            O => \N__57972\,
            I => \N__57443\
        );

    \I__14493\ : ClkMux
    port map (
            O => \N__57971\,
            I => \N__57443\
        );

    \I__14492\ : ClkMux
    port map (
            O => \N__57970\,
            I => \N__57443\
        );

    \I__14491\ : ClkMux
    port map (
            O => \N__57969\,
            I => \N__57443\
        );

    \I__14490\ : ClkMux
    port map (
            O => \N__57968\,
            I => \N__57443\
        );

    \I__14489\ : ClkMux
    port map (
            O => \N__57967\,
            I => \N__57443\
        );

    \I__14488\ : ClkMux
    port map (
            O => \N__57966\,
            I => \N__57443\
        );

    \I__14487\ : ClkMux
    port map (
            O => \N__57965\,
            I => \N__57443\
        );

    \I__14486\ : ClkMux
    port map (
            O => \N__57964\,
            I => \N__57443\
        );

    \I__14485\ : ClkMux
    port map (
            O => \N__57963\,
            I => \N__57443\
        );

    \I__14484\ : ClkMux
    port map (
            O => \N__57962\,
            I => \N__57443\
        );

    \I__14483\ : ClkMux
    port map (
            O => \N__57961\,
            I => \N__57443\
        );

    \I__14482\ : ClkMux
    port map (
            O => \N__57960\,
            I => \N__57443\
        );

    \I__14481\ : ClkMux
    port map (
            O => \N__57959\,
            I => \N__57443\
        );

    \I__14480\ : ClkMux
    port map (
            O => \N__57958\,
            I => \N__57443\
        );

    \I__14479\ : ClkMux
    port map (
            O => \N__57957\,
            I => \N__57443\
        );

    \I__14478\ : ClkMux
    port map (
            O => \N__57956\,
            I => \N__57443\
        );

    \I__14477\ : ClkMux
    port map (
            O => \N__57955\,
            I => \N__57443\
        );

    \I__14476\ : ClkMux
    port map (
            O => \N__57954\,
            I => \N__57443\
        );

    \I__14475\ : ClkMux
    port map (
            O => \N__57953\,
            I => \N__57443\
        );

    \I__14474\ : ClkMux
    port map (
            O => \N__57952\,
            I => \N__57443\
        );

    \I__14473\ : ClkMux
    port map (
            O => \N__57951\,
            I => \N__57443\
        );

    \I__14472\ : ClkMux
    port map (
            O => \N__57950\,
            I => \N__57443\
        );

    \I__14471\ : ClkMux
    port map (
            O => \N__57949\,
            I => \N__57443\
        );

    \I__14470\ : ClkMux
    port map (
            O => \N__57948\,
            I => \N__57443\
        );

    \I__14469\ : ClkMux
    port map (
            O => \N__57947\,
            I => \N__57443\
        );

    \I__14468\ : ClkMux
    port map (
            O => \N__57946\,
            I => \N__57443\
        );

    \I__14467\ : ClkMux
    port map (
            O => \N__57945\,
            I => \N__57443\
        );

    \I__14466\ : ClkMux
    port map (
            O => \N__57944\,
            I => \N__57443\
        );

    \I__14465\ : ClkMux
    port map (
            O => \N__57943\,
            I => \N__57443\
        );

    \I__14464\ : ClkMux
    port map (
            O => \N__57942\,
            I => \N__57443\
        );

    \I__14463\ : ClkMux
    port map (
            O => \N__57941\,
            I => \N__57443\
        );

    \I__14462\ : ClkMux
    port map (
            O => \N__57940\,
            I => \N__57443\
        );

    \I__14461\ : ClkMux
    port map (
            O => \N__57939\,
            I => \N__57443\
        );

    \I__14460\ : ClkMux
    port map (
            O => \N__57938\,
            I => \N__57443\
        );

    \I__14459\ : ClkMux
    port map (
            O => \N__57937\,
            I => \N__57443\
        );

    \I__14458\ : ClkMux
    port map (
            O => \N__57936\,
            I => \N__57443\
        );

    \I__14457\ : ClkMux
    port map (
            O => \N__57935\,
            I => \N__57443\
        );

    \I__14456\ : ClkMux
    port map (
            O => \N__57934\,
            I => \N__57443\
        );

    \I__14455\ : ClkMux
    port map (
            O => \N__57933\,
            I => \N__57443\
        );

    \I__14454\ : ClkMux
    port map (
            O => \N__57932\,
            I => \N__57443\
        );

    \I__14453\ : ClkMux
    port map (
            O => \N__57931\,
            I => \N__57443\
        );

    \I__14452\ : ClkMux
    port map (
            O => \N__57930\,
            I => \N__57443\
        );

    \I__14451\ : ClkMux
    port map (
            O => \N__57929\,
            I => \N__57443\
        );

    \I__14450\ : ClkMux
    port map (
            O => \N__57928\,
            I => \N__57443\
        );

    \I__14449\ : ClkMux
    port map (
            O => \N__57927\,
            I => \N__57443\
        );

    \I__14448\ : ClkMux
    port map (
            O => \N__57926\,
            I => \N__57443\
        );

    \I__14447\ : ClkMux
    port map (
            O => \N__57925\,
            I => \N__57443\
        );

    \I__14446\ : ClkMux
    port map (
            O => \N__57924\,
            I => \N__57443\
        );

    \I__14445\ : ClkMux
    port map (
            O => \N__57923\,
            I => \N__57443\
        );

    \I__14444\ : ClkMux
    port map (
            O => \N__57922\,
            I => \N__57443\
        );

    \I__14443\ : ClkMux
    port map (
            O => \N__57921\,
            I => \N__57443\
        );

    \I__14442\ : ClkMux
    port map (
            O => \N__57920\,
            I => \N__57443\
        );

    \I__14441\ : ClkMux
    port map (
            O => \N__57919\,
            I => \N__57443\
        );

    \I__14440\ : ClkMux
    port map (
            O => \N__57918\,
            I => \N__57443\
        );

    \I__14439\ : ClkMux
    port map (
            O => \N__57917\,
            I => \N__57443\
        );

    \I__14438\ : ClkMux
    port map (
            O => \N__57916\,
            I => \N__57443\
        );

    \I__14437\ : ClkMux
    port map (
            O => \N__57915\,
            I => \N__57443\
        );

    \I__14436\ : ClkMux
    port map (
            O => \N__57914\,
            I => \N__57443\
        );

    \I__14435\ : ClkMux
    port map (
            O => \N__57913\,
            I => \N__57443\
        );

    \I__14434\ : ClkMux
    port map (
            O => \N__57912\,
            I => \N__57443\
        );

    \I__14433\ : ClkMux
    port map (
            O => \N__57911\,
            I => \N__57443\
        );

    \I__14432\ : ClkMux
    port map (
            O => \N__57910\,
            I => \N__57443\
        );

    \I__14431\ : ClkMux
    port map (
            O => \N__57909\,
            I => \N__57443\
        );

    \I__14430\ : ClkMux
    port map (
            O => \N__57908\,
            I => \N__57443\
        );

    \I__14429\ : ClkMux
    port map (
            O => \N__57907\,
            I => \N__57443\
        );

    \I__14428\ : ClkMux
    port map (
            O => \N__57906\,
            I => \N__57443\
        );

    \I__14427\ : ClkMux
    port map (
            O => \N__57905\,
            I => \N__57443\
        );

    \I__14426\ : ClkMux
    port map (
            O => \N__57904\,
            I => \N__57443\
        );

    \I__14425\ : ClkMux
    port map (
            O => \N__57903\,
            I => \N__57443\
        );

    \I__14424\ : ClkMux
    port map (
            O => \N__57902\,
            I => \N__57443\
        );

    \I__14423\ : ClkMux
    port map (
            O => \N__57901\,
            I => \N__57443\
        );

    \I__14422\ : ClkMux
    port map (
            O => \N__57900\,
            I => \N__57443\
        );

    \I__14421\ : ClkMux
    port map (
            O => \N__57899\,
            I => \N__57443\
        );

    \I__14420\ : ClkMux
    port map (
            O => \N__57898\,
            I => \N__57443\
        );

    \I__14419\ : ClkMux
    port map (
            O => \N__57897\,
            I => \N__57443\
        );

    \I__14418\ : ClkMux
    port map (
            O => \N__57896\,
            I => \N__57443\
        );

    \I__14417\ : ClkMux
    port map (
            O => \N__57895\,
            I => \N__57443\
        );

    \I__14416\ : ClkMux
    port map (
            O => \N__57894\,
            I => \N__57443\
        );

    \I__14415\ : ClkMux
    port map (
            O => \N__57893\,
            I => \N__57443\
        );

    \I__14414\ : ClkMux
    port map (
            O => \N__57892\,
            I => \N__57443\
        );

    \I__14413\ : ClkMux
    port map (
            O => \N__57891\,
            I => \N__57443\
        );

    \I__14412\ : ClkMux
    port map (
            O => \N__57890\,
            I => \N__57443\
        );

    \I__14411\ : ClkMux
    port map (
            O => \N__57889\,
            I => \N__57443\
        );

    \I__14410\ : ClkMux
    port map (
            O => \N__57888\,
            I => \N__57443\
        );

    \I__14409\ : ClkMux
    port map (
            O => \N__57887\,
            I => \N__57443\
        );

    \I__14408\ : ClkMux
    port map (
            O => \N__57886\,
            I => \N__57443\
        );

    \I__14407\ : ClkMux
    port map (
            O => \N__57885\,
            I => \N__57443\
        );

    \I__14406\ : ClkMux
    port map (
            O => \N__57884\,
            I => \N__57443\
        );

    \I__14405\ : ClkMux
    port map (
            O => \N__57883\,
            I => \N__57443\
        );

    \I__14404\ : ClkMux
    port map (
            O => \N__57882\,
            I => \N__57443\
        );

    \I__14403\ : ClkMux
    port map (
            O => \N__57881\,
            I => \N__57443\
        );

    \I__14402\ : ClkMux
    port map (
            O => \N__57880\,
            I => \N__57443\
        );

    \I__14401\ : ClkMux
    port map (
            O => \N__57879\,
            I => \N__57443\
        );

    \I__14400\ : ClkMux
    port map (
            O => \N__57878\,
            I => \N__57443\
        );

    \I__14399\ : ClkMux
    port map (
            O => \N__57877\,
            I => \N__57443\
        );

    \I__14398\ : ClkMux
    port map (
            O => \N__57876\,
            I => \N__57443\
        );

    \I__14397\ : ClkMux
    port map (
            O => \N__57875\,
            I => \N__57443\
        );

    \I__14396\ : ClkMux
    port map (
            O => \N__57874\,
            I => \N__57443\
        );

    \I__14395\ : ClkMux
    port map (
            O => \N__57873\,
            I => \N__57443\
        );

    \I__14394\ : ClkMux
    port map (
            O => \N__57872\,
            I => \N__57443\
        );

    \I__14393\ : ClkMux
    port map (
            O => \N__57871\,
            I => \N__57443\
        );

    \I__14392\ : ClkMux
    port map (
            O => \N__57870\,
            I => \N__57443\
        );

    \I__14391\ : ClkMux
    port map (
            O => \N__57869\,
            I => \N__57443\
        );

    \I__14390\ : ClkMux
    port map (
            O => \N__57868\,
            I => \N__57443\
        );

    \I__14389\ : ClkMux
    port map (
            O => \N__57867\,
            I => \N__57443\
        );

    \I__14388\ : ClkMux
    port map (
            O => \N__57866\,
            I => \N__57443\
        );

    \I__14387\ : ClkMux
    port map (
            O => \N__57865\,
            I => \N__57443\
        );

    \I__14386\ : ClkMux
    port map (
            O => \N__57864\,
            I => \N__57443\
        );

    \I__14385\ : ClkMux
    port map (
            O => \N__57863\,
            I => \N__57443\
        );

    \I__14384\ : ClkMux
    port map (
            O => \N__57862\,
            I => \N__57443\
        );

    \I__14383\ : ClkMux
    port map (
            O => \N__57861\,
            I => \N__57443\
        );

    \I__14382\ : ClkMux
    port map (
            O => \N__57860\,
            I => \N__57443\
        );

    \I__14381\ : ClkMux
    port map (
            O => \N__57859\,
            I => \N__57443\
        );

    \I__14380\ : ClkMux
    port map (
            O => \N__57858\,
            I => \N__57443\
        );

    \I__14379\ : ClkMux
    port map (
            O => \N__57857\,
            I => \N__57443\
        );

    \I__14378\ : ClkMux
    port map (
            O => \N__57856\,
            I => \N__57443\
        );

    \I__14377\ : ClkMux
    port map (
            O => \N__57855\,
            I => \N__57443\
        );

    \I__14376\ : ClkMux
    port map (
            O => \N__57854\,
            I => \N__57443\
        );

    \I__14375\ : ClkMux
    port map (
            O => \N__57853\,
            I => \N__57443\
        );

    \I__14374\ : ClkMux
    port map (
            O => \N__57852\,
            I => \N__57443\
        );

    \I__14373\ : ClkMux
    port map (
            O => \N__57851\,
            I => \N__57443\
        );

    \I__14372\ : ClkMux
    port map (
            O => \N__57850\,
            I => \N__57443\
        );

    \I__14371\ : ClkMux
    port map (
            O => \N__57849\,
            I => \N__57443\
        );

    \I__14370\ : ClkMux
    port map (
            O => \N__57848\,
            I => \N__57443\
        );

    \I__14369\ : ClkMux
    port map (
            O => \N__57847\,
            I => \N__57443\
        );

    \I__14368\ : ClkMux
    port map (
            O => \N__57846\,
            I => \N__57443\
        );

    \I__14367\ : ClkMux
    port map (
            O => \N__57845\,
            I => \N__57443\
        );

    \I__14366\ : ClkMux
    port map (
            O => \N__57844\,
            I => \N__57443\
        );

    \I__14365\ : ClkMux
    port map (
            O => \N__57843\,
            I => \N__57443\
        );

    \I__14364\ : ClkMux
    port map (
            O => \N__57842\,
            I => \N__57443\
        );

    \I__14363\ : ClkMux
    port map (
            O => \N__57841\,
            I => \N__57443\
        );

    \I__14362\ : ClkMux
    port map (
            O => \N__57840\,
            I => \N__57443\
        );

    \I__14361\ : ClkMux
    port map (
            O => \N__57839\,
            I => \N__57443\
        );

    \I__14360\ : ClkMux
    port map (
            O => \N__57838\,
            I => \N__57443\
        );

    \I__14359\ : ClkMux
    port map (
            O => \N__57837\,
            I => \N__57443\
        );

    \I__14358\ : ClkMux
    port map (
            O => \N__57836\,
            I => \N__57443\
        );

    \I__14357\ : ClkMux
    port map (
            O => \N__57835\,
            I => \N__57443\
        );

    \I__14356\ : ClkMux
    port map (
            O => \N__57834\,
            I => \N__57443\
        );

    \I__14355\ : ClkMux
    port map (
            O => \N__57833\,
            I => \N__57443\
        );

    \I__14354\ : ClkMux
    port map (
            O => \N__57832\,
            I => \N__57443\
        );

    \I__14353\ : ClkMux
    port map (
            O => \N__57831\,
            I => \N__57443\
        );

    \I__14352\ : ClkMux
    port map (
            O => \N__57830\,
            I => \N__57443\
        );

    \I__14351\ : ClkMux
    port map (
            O => \N__57829\,
            I => \N__57443\
        );

    \I__14350\ : ClkMux
    port map (
            O => \N__57828\,
            I => \N__57443\
        );

    \I__14349\ : ClkMux
    port map (
            O => \N__57827\,
            I => \N__57443\
        );

    \I__14348\ : ClkMux
    port map (
            O => \N__57826\,
            I => \N__57443\
        );

    \I__14347\ : ClkMux
    port map (
            O => \N__57825\,
            I => \N__57443\
        );

    \I__14346\ : ClkMux
    port map (
            O => \N__57824\,
            I => \N__57443\
        );

    \I__14345\ : ClkMux
    port map (
            O => \N__57823\,
            I => \N__57443\
        );

    \I__14344\ : ClkMux
    port map (
            O => \N__57822\,
            I => \N__57443\
        );

    \I__14343\ : ClkMux
    port map (
            O => \N__57821\,
            I => \N__57443\
        );

    \I__14342\ : ClkMux
    port map (
            O => \N__57820\,
            I => \N__57443\
        );

    \I__14341\ : ClkMux
    port map (
            O => \N__57819\,
            I => \N__57443\
        );

    \I__14340\ : ClkMux
    port map (
            O => \N__57818\,
            I => \N__57443\
        );

    \I__14339\ : ClkMux
    port map (
            O => \N__57817\,
            I => \N__57443\
        );

    \I__14338\ : ClkMux
    port map (
            O => \N__57816\,
            I => \N__57443\
        );

    \I__14337\ : ClkMux
    port map (
            O => \N__57815\,
            I => \N__57443\
        );

    \I__14336\ : ClkMux
    port map (
            O => \N__57814\,
            I => \N__57443\
        );

    \I__14335\ : ClkMux
    port map (
            O => \N__57813\,
            I => \N__57443\
        );

    \I__14334\ : ClkMux
    port map (
            O => \N__57812\,
            I => \N__57443\
        );

    \I__14333\ : ClkMux
    port map (
            O => \N__57811\,
            I => \N__57443\
        );

    \I__14332\ : ClkMux
    port map (
            O => \N__57810\,
            I => \N__57443\
        );

    \I__14331\ : ClkMux
    port map (
            O => \N__57809\,
            I => \N__57443\
        );

    \I__14330\ : ClkMux
    port map (
            O => \N__57808\,
            I => \N__57443\
        );

    \I__14329\ : ClkMux
    port map (
            O => \N__57807\,
            I => \N__57443\
        );

    \I__14328\ : ClkMux
    port map (
            O => \N__57806\,
            I => \N__57443\
        );

    \I__14327\ : ClkMux
    port map (
            O => \N__57805\,
            I => \N__57443\
        );

    \I__14326\ : ClkMux
    port map (
            O => \N__57804\,
            I => \N__57443\
        );

    \I__14325\ : GlobalMux
    port map (
            O => \N__57443\,
            I => \clk_32MHz\
        );

    \I__14324\ : SRMux
    port map (
            O => \N__57440\,
            I => \N__57437\
        );

    \I__14323\ : LocalMux
    port map (
            O => \N__57437\,
            I => \N__57434\
        );

    \I__14322\ : Span4Mux_h
    port map (
            O => \N__57434\,
            I => \N__57431\
        );

    \I__14321\ : Span4Mux_v
    port map (
            O => \N__57431\,
            I => \N__57428\
        );

    \I__14320\ : Odrv4
    port map (
            O => \N__57428\,
            I => \comm_spi.iclk_N_764\
        );

    \I__14319\ : CascadeMux
    port map (
            O => \N__57425\,
            I => \N__57419\
        );

    \I__14318\ : CascadeMux
    port map (
            O => \N__57424\,
            I => \N__57415\
        );

    \I__14317\ : CascadeMux
    port map (
            O => \N__57423\,
            I => \N__57411\
        );

    \I__14316\ : InMux
    port map (
            O => \N__57422\,
            I => \N__57395\
        );

    \I__14315\ : InMux
    port map (
            O => \N__57419\,
            I => \N__57395\
        );

    \I__14314\ : InMux
    port map (
            O => \N__57418\,
            I => \N__57395\
        );

    \I__14313\ : InMux
    port map (
            O => \N__57415\,
            I => \N__57395\
        );

    \I__14312\ : InMux
    port map (
            O => \N__57414\,
            I => \N__57395\
        );

    \I__14311\ : InMux
    port map (
            O => \N__57411\,
            I => \N__57395\
        );

    \I__14310\ : InMux
    port map (
            O => \N__57410\,
            I => \N__57395\
        );

    \I__14309\ : LocalMux
    port map (
            O => \N__57395\,
            I => \N__57385\
        );

    \I__14308\ : CascadeMux
    port map (
            O => \N__57394\,
            I => \N__57376\
        );

    \I__14307\ : CascadeMux
    port map (
            O => \N__57393\,
            I => \N__57370\
        );

    \I__14306\ : CascadeMux
    port map (
            O => \N__57392\,
            I => \N__57366\
        );

    \I__14305\ : CascadeMux
    port map (
            O => \N__57391\,
            I => \N__57362\
        );

    \I__14304\ : CascadeMux
    port map (
            O => \N__57390\,
            I => \N__57358\
        );

    \I__14303\ : CascadeMux
    port map (
            O => \N__57389\,
            I => \N__57354\
        );

    \I__14302\ : CascadeMux
    port map (
            O => \N__57388\,
            I => \N__57350\
        );

    \I__14301\ : Span4Mux_v
    port map (
            O => \N__57385\,
            I => \N__57347\
        );

    \I__14300\ : CascadeMux
    port map (
            O => \N__57384\,
            I => \N__57343\
        );

    \I__14299\ : CascadeMux
    port map (
            O => \N__57383\,
            I => \N__57339\
        );

    \I__14298\ : CascadeMux
    port map (
            O => \N__57382\,
            I => \N__57335\
        );

    \I__14297\ : CascadeMux
    port map (
            O => \N__57381\,
            I => \N__57331\
        );

    \I__14296\ : SRMux
    port map (
            O => \N__57380\,
            I => \N__57328\
        );

    \I__14295\ : SRMux
    port map (
            O => \N__57379\,
            I => \N__57321\
        );

    \I__14294\ : InMux
    port map (
            O => \N__57376\,
            I => \N__57301\
        );

    \I__14293\ : InMux
    port map (
            O => \N__57375\,
            I => \N__57301\
        );

    \I__14292\ : InMux
    port map (
            O => \N__57374\,
            I => \N__57301\
        );

    \I__14291\ : InMux
    port map (
            O => \N__57373\,
            I => \N__57301\
        );

    \I__14290\ : InMux
    port map (
            O => \N__57370\,
            I => \N__57301\
        );

    \I__14289\ : InMux
    port map (
            O => \N__57369\,
            I => \N__57301\
        );

    \I__14288\ : InMux
    port map (
            O => \N__57366\,
            I => \N__57301\
        );

    \I__14287\ : InMux
    port map (
            O => \N__57365\,
            I => \N__57301\
        );

    \I__14286\ : InMux
    port map (
            O => \N__57362\,
            I => \N__57286\
        );

    \I__14285\ : InMux
    port map (
            O => \N__57361\,
            I => \N__57286\
        );

    \I__14284\ : InMux
    port map (
            O => \N__57358\,
            I => \N__57286\
        );

    \I__14283\ : InMux
    port map (
            O => \N__57357\,
            I => \N__57286\
        );

    \I__14282\ : InMux
    port map (
            O => \N__57354\,
            I => \N__57286\
        );

    \I__14281\ : InMux
    port map (
            O => \N__57353\,
            I => \N__57286\
        );

    \I__14280\ : InMux
    port map (
            O => \N__57350\,
            I => \N__57286\
        );

    \I__14279\ : Span4Mux_v
    port map (
            O => \N__57347\,
            I => \N__57283\
        );

    \I__14278\ : InMux
    port map (
            O => \N__57346\,
            I => \N__57266\
        );

    \I__14277\ : InMux
    port map (
            O => \N__57343\,
            I => \N__57266\
        );

    \I__14276\ : InMux
    port map (
            O => \N__57342\,
            I => \N__57266\
        );

    \I__14275\ : InMux
    port map (
            O => \N__57339\,
            I => \N__57266\
        );

    \I__14274\ : InMux
    port map (
            O => \N__57338\,
            I => \N__57266\
        );

    \I__14273\ : InMux
    port map (
            O => \N__57335\,
            I => \N__57266\
        );

    \I__14272\ : InMux
    port map (
            O => \N__57334\,
            I => \N__57266\
        );

    \I__14271\ : InMux
    port map (
            O => \N__57331\,
            I => \N__57266\
        );

    \I__14270\ : LocalMux
    port map (
            O => \N__57328\,
            I => \N__57263\
        );

    \I__14269\ : CascadeMux
    port map (
            O => \N__57327\,
            I => \N__57260\
        );

    \I__14268\ : CascadeMux
    port map (
            O => \N__57326\,
            I => \N__57256\
        );

    \I__14267\ : CascadeMux
    port map (
            O => \N__57325\,
            I => \N__57252\
        );

    \I__14266\ : CascadeMux
    port map (
            O => \N__57324\,
            I => \N__57248\
        );

    \I__14265\ : LocalMux
    port map (
            O => \N__57321\,
            I => \N__57245\
        );

    \I__14264\ : SRMux
    port map (
            O => \N__57320\,
            I => \N__57242\
        );

    \I__14263\ : SRMux
    port map (
            O => \N__57319\,
            I => \N__57239\
        );

    \I__14262\ : SRMux
    port map (
            O => \N__57318\,
            I => \N__57233\
        );

    \I__14261\ : LocalMux
    port map (
            O => \N__57301\,
            I => \N__57227\
        );

    \I__14260\ : LocalMux
    port map (
            O => \N__57286\,
            I => \N__57227\
        );

    \I__14259\ : Span4Mux_v
    port map (
            O => \N__57283\,
            I => \N__57222\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__57266\,
            I => \N__57222\
        );

    \I__14257\ : Span4Mux_h
    port map (
            O => \N__57263\,
            I => \N__57219\
        );

    \I__14256\ : InMux
    port map (
            O => \N__57260\,
            I => \N__57204\
        );

    \I__14255\ : InMux
    port map (
            O => \N__57259\,
            I => \N__57204\
        );

    \I__14254\ : InMux
    port map (
            O => \N__57256\,
            I => \N__57204\
        );

    \I__14253\ : InMux
    port map (
            O => \N__57255\,
            I => \N__57204\
        );

    \I__14252\ : InMux
    port map (
            O => \N__57252\,
            I => \N__57204\
        );

    \I__14251\ : InMux
    port map (
            O => \N__57251\,
            I => \N__57204\
        );

    \I__14250\ : InMux
    port map (
            O => \N__57248\,
            I => \N__57204\
        );

    \I__14249\ : Span4Mux_v
    port map (
            O => \N__57245\,
            I => \N__57197\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__57242\,
            I => \N__57197\
        );

    \I__14247\ : LocalMux
    port map (
            O => \N__57239\,
            I => \N__57197\
        );

    \I__14246\ : SRMux
    port map (
            O => \N__57238\,
            I => \N__57194\
        );

    \I__14245\ : InMux
    port map (
            O => \N__57237\,
            I => \N__57191\
        );

    \I__14244\ : SRMux
    port map (
            O => \N__57236\,
            I => \N__57188\
        );

    \I__14243\ : LocalMux
    port map (
            O => \N__57233\,
            I => \N__57182\
        );

    \I__14242\ : IoInMux
    port map (
            O => \N__57232\,
            I => \N__57179\
        );

    \I__14241\ : Span4Mux_v
    port map (
            O => \N__57227\,
            I => \N__57174\
        );

    \I__14240\ : Span4Mux_v
    port map (
            O => \N__57222\,
            I => \N__57174\
        );

    \I__14239\ : Span4Mux_h
    port map (
            O => \N__57219\,
            I => \N__57171\
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__57204\,
            I => \N__57168\
        );

    \I__14237\ : Span4Mux_v
    port map (
            O => \N__57197\,
            I => \N__57158\
        );

    \I__14236\ : LocalMux
    port map (
            O => \N__57194\,
            I => \N__57158\
        );

    \I__14235\ : LocalMux
    port map (
            O => \N__57191\,
            I => \N__57158\
        );

    \I__14234\ : LocalMux
    port map (
            O => \N__57188\,
            I => \N__57158\
        );

    \I__14233\ : SRMux
    port map (
            O => \N__57187\,
            I => \N__57155\
        );

    \I__14232\ : InMux
    port map (
            O => \N__57186\,
            I => \N__57152\
        );

    \I__14231\ : SRMux
    port map (
            O => \N__57185\,
            I => \N__57149\
        );

    \I__14230\ : Span12Mux_h
    port map (
            O => \N__57182\,
            I => \N__57144\
        );

    \I__14229\ : LocalMux
    port map (
            O => \N__57179\,
            I => \N__57141\
        );

    \I__14228\ : Span4Mux_h
    port map (
            O => \N__57174\,
            I => \N__57138\
        );

    \I__14227\ : Span4Mux_h
    port map (
            O => \N__57171\,
            I => \N__57133\
        );

    \I__14226\ : Span4Mux_h
    port map (
            O => \N__57168\,
            I => \N__57133\
        );

    \I__14225\ : SRMux
    port map (
            O => \N__57167\,
            I => \N__57130\
        );

    \I__14224\ : Span4Mux_v
    port map (
            O => \N__57158\,
            I => \N__57121\
        );

    \I__14223\ : LocalMux
    port map (
            O => \N__57155\,
            I => \N__57121\
        );

    \I__14222\ : LocalMux
    port map (
            O => \N__57152\,
            I => \N__57121\
        );

    \I__14221\ : LocalMux
    port map (
            O => \N__57149\,
            I => \N__57121\
        );

    \I__14220\ : SRMux
    port map (
            O => \N__57148\,
            I => \N__57118\
        );

    \I__14219\ : SRMux
    port map (
            O => \N__57147\,
            I => \N__57115\
        );

    \I__14218\ : Span12Mux_h
    port map (
            O => \N__57144\,
            I => \N__57112\
        );

    \I__14217\ : Span12Mux_s8_v
    port map (
            O => \N__57141\,
            I => \N__57109\
        );

    \I__14216\ : Span4Mux_h
    port map (
            O => \N__57138\,
            I => \N__57106\
        );

    \I__14215\ : Span4Mux_h
    port map (
            O => \N__57133\,
            I => \N__57103\
        );

    \I__14214\ : LocalMux
    port map (
            O => \N__57130\,
            I => \N__57100\
        );

    \I__14213\ : Span4Mux_v
    port map (
            O => \N__57121\,
            I => \N__57093\
        );

    \I__14212\ : LocalMux
    port map (
            O => \N__57118\,
            I => \N__57093\
        );

    \I__14211\ : LocalMux
    port map (
            O => \N__57115\,
            I => \N__57093\
        );

    \I__14210\ : Odrv12
    port map (
            O => \N__57112\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14209\ : Odrv12
    port map (
            O => \N__57109\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14208\ : Odrv4
    port map (
            O => \N__57106\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14207\ : Odrv4
    port map (
            O => \N__57103\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14206\ : Odrv4
    port map (
            O => \N__57100\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14205\ : Odrv4
    port map (
            O => \N__57093\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14204\ : InMux
    port map (
            O => \N__57080\,
            I => \N__57076\
        );

    \I__14203\ : InMux
    port map (
            O => \N__57079\,
            I => \N__57073\
        );

    \I__14202\ : LocalMux
    port map (
            O => \N__57076\,
            I => \N__57070\
        );

    \I__14201\ : LocalMux
    port map (
            O => \N__57073\,
            I => \N__57067\
        );

    \I__14200\ : Odrv12
    port map (
            O => \N__57070\,
            I => \comm_spi.n14609\
        );

    \I__14199\ : Odrv4
    port map (
            O => \N__57067\,
            I => \comm_spi.n14609\
        );

    \I__14198\ : ClkMux
    port map (
            O => \N__57062\,
            I => \N__57059\
        );

    \I__14197\ : LocalMux
    port map (
            O => \N__57059\,
            I => \N__57055\
        );

    \I__14196\ : ClkMux
    port map (
            O => \N__57058\,
            I => \N__57052\
        );

    \I__14195\ : Span4Mux_h
    port map (
            O => \N__57055\,
            I => \N__57044\
        );

    \I__14194\ : LocalMux
    port map (
            O => \N__57052\,
            I => \N__57044\
        );

    \I__14193\ : ClkMux
    port map (
            O => \N__57051\,
            I => \N__57041\
        );

    \I__14192\ : ClkMux
    port map (
            O => \N__57050\,
            I => \N__57037\
        );

    \I__14191\ : ClkMux
    port map (
            O => \N__57049\,
            I => \N__57032\
        );

    \I__14190\ : Span4Mux_v
    port map (
            O => \N__57044\,
            I => \N__57027\
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__57041\,
            I => \N__57027\
        );

    \I__14188\ : ClkMux
    port map (
            O => \N__57040\,
            I => \N__57024\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__57037\,
            I => \N__57021\
        );

    \I__14186\ : ClkMux
    port map (
            O => \N__57036\,
            I => \N__57018\
        );

    \I__14185\ : ClkMux
    port map (
            O => \N__57035\,
            I => \N__57013\
        );

    \I__14184\ : LocalMux
    port map (
            O => \N__57032\,
            I => \N__57009\
        );

    \I__14183\ : Span4Mux_h
    port map (
            O => \N__57027\,
            I => \N__57004\
        );

    \I__14182\ : LocalMux
    port map (
            O => \N__57024\,
            I => \N__57004\
        );

    \I__14181\ : Span4Mux_v
    port map (
            O => \N__57021\,
            I => \N__56999\
        );

    \I__14180\ : LocalMux
    port map (
            O => \N__57018\,
            I => \N__56999\
        );

    \I__14179\ : ClkMux
    port map (
            O => \N__57017\,
            I => \N__56992\
        );

    \I__14178\ : ClkMux
    port map (
            O => \N__57016\,
            I => \N__56988\
        );

    \I__14177\ : LocalMux
    port map (
            O => \N__57013\,
            I => \N__56984\
        );

    \I__14176\ : ClkMux
    port map (
            O => \N__57012\,
            I => \N__56980\
        );

    \I__14175\ : Span4Mux_v
    port map (
            O => \N__57009\,
            I => \N__56975\
        );

    \I__14174\ : Span4Mux_v
    port map (
            O => \N__57004\,
            I => \N__56975\
        );

    \I__14173\ : Span4Mux_h
    port map (
            O => \N__56999\,
            I => \N__56972\
        );

    \I__14172\ : ClkMux
    port map (
            O => \N__56998\,
            I => \N__56969\
        );

    \I__14171\ : ClkMux
    port map (
            O => \N__56997\,
            I => \N__56966\
        );

    \I__14170\ : ClkMux
    port map (
            O => \N__56996\,
            I => \N__56963\
        );

    \I__14169\ : ClkMux
    port map (
            O => \N__56995\,
            I => \N__56960\
        );

    \I__14168\ : LocalMux
    port map (
            O => \N__56992\,
            I => \N__56957\
        );

    \I__14167\ : ClkMux
    port map (
            O => \N__56991\,
            I => \N__56954\
        );

    \I__14166\ : LocalMux
    port map (
            O => \N__56988\,
            I => \N__56951\
        );

    \I__14165\ : ClkMux
    port map (
            O => \N__56987\,
            I => \N__56948\
        );

    \I__14164\ : Span4Mux_v
    port map (
            O => \N__56984\,
            I => \N__56945\
        );

    \I__14163\ : ClkMux
    port map (
            O => \N__56983\,
            I => \N__56942\
        );

    \I__14162\ : LocalMux
    port map (
            O => \N__56980\,
            I => \N__56939\
        );

    \I__14161\ : Span4Mux_h
    port map (
            O => \N__56975\,
            I => \N__56936\
        );

    \I__14160\ : Span4Mux_v
    port map (
            O => \N__56972\,
            I => \N__56931\
        );

    \I__14159\ : LocalMux
    port map (
            O => \N__56969\,
            I => \N__56931\
        );

    \I__14158\ : LocalMux
    port map (
            O => \N__56966\,
            I => \N__56926\
        );

    \I__14157\ : LocalMux
    port map (
            O => \N__56963\,
            I => \N__56926\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__56960\,
            I => \N__56919\
        );

    \I__14155\ : Span4Mux_h
    port map (
            O => \N__56957\,
            I => \N__56919\
        );

    \I__14154\ : LocalMux
    port map (
            O => \N__56954\,
            I => \N__56919\
        );

    \I__14153\ : Span4Mux_h
    port map (
            O => \N__56951\,
            I => \N__56912\
        );

    \I__14152\ : LocalMux
    port map (
            O => \N__56948\,
            I => \N__56912\
        );

    \I__14151\ : Span4Mux_h
    port map (
            O => \N__56945\,
            I => \N__56907\
        );

    \I__14150\ : LocalMux
    port map (
            O => \N__56942\,
            I => \N__56904\
        );

    \I__14149\ : Span4Mux_v
    port map (
            O => \N__56939\,
            I => \N__56899\
        );

    \I__14148\ : Span4Mux_v
    port map (
            O => \N__56936\,
            I => \N__56899\
        );

    \I__14147\ : Span4Mux_v
    port map (
            O => \N__56931\,
            I => \N__56892\
        );

    \I__14146\ : Span4Mux_v
    port map (
            O => \N__56926\,
            I => \N__56892\
        );

    \I__14145\ : Span4Mux_v
    port map (
            O => \N__56919\,
            I => \N__56892\
        );

    \I__14144\ : ClkMux
    port map (
            O => \N__56918\,
            I => \N__56889\
        );

    \I__14143\ : ClkMux
    port map (
            O => \N__56917\,
            I => \N__56886\
        );

    \I__14142\ : Span4Mux_v
    port map (
            O => \N__56912\,
            I => \N__56883\
        );

    \I__14141\ : ClkMux
    port map (
            O => \N__56911\,
            I => \N__56880\
        );

    \I__14140\ : ClkMux
    port map (
            O => \N__56910\,
            I => \N__56877\
        );

    \I__14139\ : Odrv4
    port map (
            O => \N__56907\,
            I => \comm_spi.iclk\
        );

    \I__14138\ : Odrv12
    port map (
            O => \N__56904\,
            I => \comm_spi.iclk\
        );

    \I__14137\ : Odrv4
    port map (
            O => \N__56899\,
            I => \comm_spi.iclk\
        );

    \I__14136\ : Odrv4
    port map (
            O => \N__56892\,
            I => \comm_spi.iclk\
        );

    \I__14135\ : LocalMux
    port map (
            O => \N__56889\,
            I => \comm_spi.iclk\
        );

    \I__14134\ : LocalMux
    port map (
            O => \N__56886\,
            I => \comm_spi.iclk\
        );

    \I__14133\ : Odrv4
    port map (
            O => \N__56883\,
            I => \comm_spi.iclk\
        );

    \I__14132\ : LocalMux
    port map (
            O => \N__56880\,
            I => \comm_spi.iclk\
        );

    \I__14131\ : LocalMux
    port map (
            O => \N__56877\,
            I => \comm_spi.iclk\
        );

    \I__14130\ : SRMux
    port map (
            O => \N__56858\,
            I => \N__56855\
        );

    \I__14129\ : LocalMux
    port map (
            O => \N__56855\,
            I => \N__56849\
        );

    \I__14128\ : SRMux
    port map (
            O => \N__56854\,
            I => \N__56846\
        );

    \I__14127\ : CascadeMux
    port map (
            O => \N__56853\,
            I => \N__56838\
        );

    \I__14126\ : InMux
    port map (
            O => \N__56852\,
            I => \N__56829\
        );

    \I__14125\ : Span4Mux_v
    port map (
            O => \N__56849\,
            I => \N__56824\
        );

    \I__14124\ : LocalMux
    port map (
            O => \N__56846\,
            I => \N__56824\
        );

    \I__14123\ : InMux
    port map (
            O => \N__56845\,
            I => \N__56818\
        );

    \I__14122\ : InMux
    port map (
            O => \N__56844\,
            I => \N__56818\
        );

    \I__14121\ : InMux
    port map (
            O => \N__56843\,
            I => \N__56811\
        );

    \I__14120\ : InMux
    port map (
            O => \N__56842\,
            I => \N__56811\
        );

    \I__14119\ : InMux
    port map (
            O => \N__56841\,
            I => \N__56804\
        );

    \I__14118\ : InMux
    port map (
            O => \N__56838\,
            I => \N__56795\
        );

    \I__14117\ : InMux
    port map (
            O => \N__56837\,
            I => \N__56795\
        );

    \I__14116\ : InMux
    port map (
            O => \N__56836\,
            I => \N__56795\
        );

    \I__14115\ : InMux
    port map (
            O => \N__56835\,
            I => \N__56795\
        );

    \I__14114\ : InMux
    port map (
            O => \N__56834\,
            I => \N__56792\
        );

    \I__14113\ : InMux
    port map (
            O => \N__56833\,
            I => \N__56787\
        );

    \I__14112\ : InMux
    port map (
            O => \N__56832\,
            I => \N__56787\
        );

    \I__14111\ : LocalMux
    port map (
            O => \N__56829\,
            I => \N__56784\
        );

    \I__14110\ : Span4Mux_v
    port map (
            O => \N__56824\,
            I => \N__56781\
        );

    \I__14109\ : SRMux
    port map (
            O => \N__56823\,
            I => \N__56778\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__56818\,
            I => \N__56772\
        );

    \I__14107\ : InMux
    port map (
            O => \N__56817\,
            I => \N__56767\
        );

    \I__14106\ : InMux
    port map (
            O => \N__56816\,
            I => \N__56767\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56764\
        );

    \I__14104\ : InMux
    port map (
            O => \N__56810\,
            I => \N__56761\
        );

    \I__14103\ : InMux
    port map (
            O => \N__56809\,
            I => \N__56755\
        );

    \I__14102\ : InMux
    port map (
            O => \N__56808\,
            I => \N__56755\
        );

    \I__14101\ : InMux
    port map (
            O => \N__56807\,
            I => \N__56752\
        );

    \I__14100\ : LocalMux
    port map (
            O => \N__56804\,
            I => \N__56737\
        );

    \I__14099\ : LocalMux
    port map (
            O => \N__56795\,
            I => \N__56737\
        );

    \I__14098\ : LocalMux
    port map (
            O => \N__56792\,
            I => \N__56732\
        );

    \I__14097\ : LocalMux
    port map (
            O => \N__56787\,
            I => \N__56732\
        );

    \I__14096\ : Span4Mux_v
    port map (
            O => \N__56784\,
            I => \N__56727\
        );

    \I__14095\ : Span4Mux_v
    port map (
            O => \N__56781\,
            I => \N__56727\
        );

    \I__14094\ : LocalMux
    port map (
            O => \N__56778\,
            I => \N__56724\
        );

    \I__14093\ : InMux
    port map (
            O => \N__56777\,
            I => \N__56719\
        );

    \I__14092\ : InMux
    port map (
            O => \N__56776\,
            I => \N__56719\
        );

    \I__14091\ : InMux
    port map (
            O => \N__56775\,
            I => \N__56716\
        );

    \I__14090\ : Span4Mux_h
    port map (
            O => \N__56772\,
            I => \N__56713\
        );

    \I__14089\ : LocalMux
    port map (
            O => \N__56767\,
            I => \N__56706\
        );

    \I__14088\ : Span4Mux_v
    port map (
            O => \N__56764\,
            I => \N__56706\
        );

    \I__14087\ : LocalMux
    port map (
            O => \N__56761\,
            I => \N__56706\
        );

    \I__14086\ : InMux
    port map (
            O => \N__56760\,
            I => \N__56703\
        );

    \I__14085\ : LocalMux
    port map (
            O => \N__56755\,
            I => \N__56698\
        );

    \I__14084\ : LocalMux
    port map (
            O => \N__56752\,
            I => \N__56698\
        );

    \I__14083\ : InMux
    port map (
            O => \N__56751\,
            I => \N__56695\
        );

    \I__14082\ : InMux
    port map (
            O => \N__56750\,
            I => \N__56684\
        );

    \I__14081\ : InMux
    port map (
            O => \N__56749\,
            I => \N__56684\
        );

    \I__14080\ : InMux
    port map (
            O => \N__56748\,
            I => \N__56684\
        );

    \I__14079\ : InMux
    port map (
            O => \N__56747\,
            I => \N__56684\
        );

    \I__14078\ : InMux
    port map (
            O => \N__56746\,
            I => \N__56684\
        );

    \I__14077\ : InMux
    port map (
            O => \N__56745\,
            I => \N__56675\
        );

    \I__14076\ : InMux
    port map (
            O => \N__56744\,
            I => \N__56675\
        );

    \I__14075\ : InMux
    port map (
            O => \N__56743\,
            I => \N__56675\
        );

    \I__14074\ : InMux
    port map (
            O => \N__56742\,
            I => \N__56675\
        );

    \I__14073\ : Span4Mux_v
    port map (
            O => \N__56737\,
            I => \N__56672\
        );

    \I__14072\ : Span4Mux_h
    port map (
            O => \N__56732\,
            I => \N__56667\
        );

    \I__14071\ : Span4Mux_h
    port map (
            O => \N__56727\,
            I => \N__56667\
        );

    \I__14070\ : Span12Mux_h
    port map (
            O => \N__56724\,
            I => \N__56662\
        );

    \I__14069\ : LocalMux
    port map (
            O => \N__56719\,
            I => \N__56662\
        );

    \I__14068\ : LocalMux
    port map (
            O => \N__56716\,
            I => \N__56655\
        );

    \I__14067\ : Span4Mux_v
    port map (
            O => \N__56713\,
            I => \N__56655\
        );

    \I__14066\ : Span4Mux_h
    port map (
            O => \N__56706\,
            I => \N__56655\
        );

    \I__14065\ : LocalMux
    port map (
            O => \N__56703\,
            I => \N__56650\
        );

    \I__14064\ : Span4Mux_v
    port map (
            O => \N__56698\,
            I => \N__56650\
        );

    \I__14063\ : LocalMux
    port map (
            O => \N__56695\,
            I => comm_clear
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__56684\,
            I => comm_clear
        );

    \I__14061\ : LocalMux
    port map (
            O => \N__56675\,
            I => comm_clear
        );

    \I__14060\ : Odrv4
    port map (
            O => \N__56672\,
            I => comm_clear
        );

    \I__14059\ : Odrv4
    port map (
            O => \N__56667\,
            I => comm_clear
        );

    \I__14058\ : Odrv12
    port map (
            O => \N__56662\,
            I => comm_clear
        );

    \I__14057\ : Odrv4
    port map (
            O => \N__56655\,
            I => comm_clear
        );

    \I__14056\ : Odrv4
    port map (
            O => \N__56650\,
            I => comm_clear
        );

    \I__14055\ : InMux
    port map (
            O => \N__56633\,
            I => \N__56629\
        );

    \I__14054\ : InMux
    port map (
            O => \N__56632\,
            I => \N__56625\
        );

    \I__14053\ : LocalMux
    port map (
            O => \N__56629\,
            I => \N__56622\
        );

    \I__14052\ : InMux
    port map (
            O => \N__56628\,
            I => \N__56619\
        );

    \I__14051\ : LocalMux
    port map (
            O => \N__56625\,
            I => \N__56616\
        );

    \I__14050\ : Span4Mux_v
    port map (
            O => \N__56622\,
            I => \N__56611\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__56619\,
            I => \N__56611\
        );

    \I__14048\ : Sp12to4
    port map (
            O => \N__56616\,
            I => \N__56608\
        );

    \I__14047\ : Span4Mux_v
    port map (
            O => \N__56611\,
            I => \N__56605\
        );

    \I__14046\ : Span12Mux_v
    port map (
            O => \N__56608\,
            I => \N__56600\
        );

    \I__14045\ : Sp12to4
    port map (
            O => \N__56605\,
            I => \N__56600\
        );

    \I__14044\ : Odrv12
    port map (
            O => \N__56600\,
            I => comm_tx_buf_0
        );

    \I__14043\ : SRMux
    port map (
            O => \N__56597\,
            I => \N__56594\
        );

    \I__14042\ : LocalMux
    port map (
            O => \N__56594\,
            I => \N__56591\
        );

    \I__14041\ : Span4Mux_h
    port map (
            O => \N__56591\,
            I => \N__56588\
        );

    \I__14040\ : Odrv4
    port map (
            O => \N__56588\,
            I => \comm_spi.data_tx_7__N_796\
        );

    \I__14039\ : InMux
    port map (
            O => \N__56585\,
            I => \N__56581\
        );

    \I__14038\ : InMux
    port map (
            O => \N__56584\,
            I => \N__56578\
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__56581\,
            I => \N__56572\
        );

    \I__14036\ : LocalMux
    port map (
            O => \N__56578\,
            I => \N__56572\
        );

    \I__14035\ : InMux
    port map (
            O => \N__56577\,
            I => \N__56569\
        );

    \I__14034\ : Odrv4
    port map (
            O => \N__56572\,
            I => \comm_spi.n22661\
        );

    \I__14033\ : LocalMux
    port map (
            O => \N__56569\,
            I => \comm_spi.n22661\
        );

    \I__14032\ : InMux
    port map (
            O => \N__56564\,
            I => \N__56560\
        );

    \I__14031\ : InMux
    port map (
            O => \N__56563\,
            I => \N__56557\
        );

    \I__14030\ : LocalMux
    port map (
            O => \N__56560\,
            I => \N__56554\
        );

    \I__14029\ : LocalMux
    port map (
            O => \N__56557\,
            I => \comm_spi.n14623\
        );

    \I__14028\ : Odrv4
    port map (
            O => \N__56554\,
            I => \comm_spi.n14623\
        );

    \I__14027\ : SRMux
    port map (
            O => \N__56549\,
            I => \N__56546\
        );

    \I__14026\ : LocalMux
    port map (
            O => \N__56546\,
            I => \N__56543\
        );

    \I__14025\ : Span4Mux_v
    port map (
            O => \N__56543\,
            I => \N__56539\
        );

    \I__14024\ : SRMux
    port map (
            O => \N__56542\,
            I => \N__56536\
        );

    \I__14023\ : Span4Mux_v
    port map (
            O => \N__56539\,
            I => \N__56530\
        );

    \I__14022\ : LocalMux
    port map (
            O => \N__56536\,
            I => \N__56530\
        );

    \I__14021\ : SRMux
    port map (
            O => \N__56535\,
            I => \N__56527\
        );

    \I__14020\ : Span4Mux_h
    port map (
            O => \N__56530\,
            I => \N__56524\
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__56527\,
            I => \N__56521\
        );

    \I__14018\ : Span4Mux_v
    port map (
            O => \N__56524\,
            I => \N__56516\
        );

    \I__14017\ : Span4Mux_v
    port map (
            O => \N__56521\,
            I => \N__56516\
        );

    \I__14016\ : Odrv4
    port map (
            O => \N__56516\,
            I => \comm_spi.data_tx_7__N_767\
        );

    \I__14015\ : InMux
    port map (
            O => \N__56513\,
            I => \N__56510\
        );

    \I__14014\ : LocalMux
    port map (
            O => \N__56510\,
            I => \N__56507\
        );

    \I__14013\ : Span4Mux_h
    port map (
            O => \N__56507\,
            I => \N__56502\
        );

    \I__14012\ : InMux
    port map (
            O => \N__56506\,
            I => \N__56499\
        );

    \I__14011\ : InMux
    port map (
            O => \N__56505\,
            I => \N__56496\
        );

    \I__14010\ : Odrv4
    port map (
            O => \N__56502\,
            I => comm_tx_buf_7
        );

    \I__14009\ : LocalMux
    port map (
            O => \N__56499\,
            I => comm_tx_buf_7
        );

    \I__14008\ : LocalMux
    port map (
            O => \N__56496\,
            I => comm_tx_buf_7
        );

    \I__14007\ : SRMux
    port map (
            O => \N__56489\,
            I => \N__56484\
        );

    \I__14006\ : SRMux
    port map (
            O => \N__56488\,
            I => \N__56481\
        );

    \I__14005\ : SRMux
    port map (
            O => \N__56487\,
            I => \N__56478\
        );

    \I__14004\ : LocalMux
    port map (
            O => \N__56484\,
            I => \N__56475\
        );

    \I__14003\ : LocalMux
    port map (
            O => \N__56481\,
            I => \N__56470\
        );

    \I__14002\ : LocalMux
    port map (
            O => \N__56478\,
            I => \N__56470\
        );

    \I__14001\ : Span4Mux_v
    port map (
            O => \N__56475\,
            I => \N__56467\
        );

    \I__14000\ : Span4Mux_v
    port map (
            O => \N__56470\,
            I => \N__56464\
        );

    \I__13999\ : Odrv4
    port map (
            O => \N__56467\,
            I => \comm_spi.data_tx_7__N_775\
        );

    \I__13998\ : Odrv4
    port map (
            O => \N__56464\,
            I => \comm_spi.data_tx_7__N_775\
        );

    \I__13997\ : InMux
    port map (
            O => \N__56459\,
            I => \N__56456\
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__56456\,
            I => \N__56452\
        );

    \I__13995\ : InMux
    port map (
            O => \N__56455\,
            I => \N__56449\
        );

    \I__13994\ : Odrv4
    port map (
            O => \N__56452\,
            I => \comm_spi.n14635\
        );

    \I__13993\ : LocalMux
    port map (
            O => \N__56449\,
            I => \comm_spi.n14635\
        );

    \I__13992\ : SRMux
    port map (
            O => \N__56444\,
            I => \N__56441\
        );

    \I__13991\ : LocalMux
    port map (
            O => \N__56441\,
            I => \N__56438\
        );

    \I__13990\ : Span4Mux_v
    port map (
            O => \N__56438\,
            I => \N__56435\
        );

    \I__13989\ : Odrv4
    port map (
            O => \N__56435\,
            I => \comm_spi.data_tx_7__N_793\
        );

    \I__13988\ : InMux
    port map (
            O => \N__56432\,
            I => \N__56429\
        );

    \I__13987\ : LocalMux
    port map (
            O => \N__56429\,
            I => \N__56426\
        );

    \I__13986\ : Span4Mux_h
    port map (
            O => \N__56426\,
            I => \N__56422\
        );

    \I__13985\ : InMux
    port map (
            O => \N__56425\,
            I => \N__56419\
        );

    \I__13984\ : Odrv4
    port map (
            O => \N__56422\,
            I => \comm_spi.n22664\
        );

    \I__13983\ : LocalMux
    port map (
            O => \N__56419\,
            I => \comm_spi.n22664\
        );

    \I__13982\ : InMux
    port map (
            O => \N__56414\,
            I => \N__56411\
        );

    \I__13981\ : LocalMux
    port map (
            O => \N__56411\,
            I => \comm_spi.n14612\
        );

    \I__13980\ : SRMux
    port map (
            O => \N__56408\,
            I => \N__56405\
        );

    \I__13979\ : LocalMux
    port map (
            O => \N__56405\,
            I => \N__56402\
        );

    \I__13978\ : Sp12to4
    port map (
            O => \N__56402\,
            I => \N__56399\
        );

    \I__13977\ : Odrv12
    port map (
            O => \N__56399\,
            I => \comm_spi.iclk_N_763\
        );

    \I__13976\ : InMux
    port map (
            O => \N__56396\,
            I => \N__56391\
        );

    \I__13975\ : InMux
    port map (
            O => \N__56395\,
            I => \N__56388\
        );

    \I__13974\ : InMux
    port map (
            O => \N__56394\,
            I => \N__56385\
        );

    \I__13973\ : LocalMux
    port map (
            O => \N__56391\,
            I => \comm_spi.n22688\
        );

    \I__13972\ : LocalMux
    port map (
            O => \N__56388\,
            I => \comm_spi.n22688\
        );

    \I__13971\ : LocalMux
    port map (
            O => \N__56385\,
            I => \comm_spi.n22688\
        );

    \I__13970\ : CascadeMux
    port map (
            O => \N__56378\,
            I => \N__56374\
        );

    \I__13969\ : InMux
    port map (
            O => \N__56377\,
            I => \N__56364\
        );

    \I__13968\ : InMux
    port map (
            O => \N__56374\,
            I => \N__56348\
        );

    \I__13967\ : InMux
    port map (
            O => \N__56373\,
            I => \N__56348\
        );

    \I__13966\ : InMux
    port map (
            O => \N__56372\,
            I => \N__56348\
        );

    \I__13965\ : InMux
    port map (
            O => \N__56371\,
            I => \N__56348\
        );

    \I__13964\ : InMux
    port map (
            O => \N__56370\,
            I => \N__56345\
        );

    \I__13963\ : InMux
    port map (
            O => \N__56369\,
            I => \N__56342\
        );

    \I__13962\ : InMux
    port map (
            O => \N__56368\,
            I => \N__56326\
        );

    \I__13961\ : InMux
    port map (
            O => \N__56367\,
            I => \N__56314\
        );

    \I__13960\ : LocalMux
    port map (
            O => \N__56364\,
            I => \N__56310\
        );

    \I__13959\ : InMux
    port map (
            O => \N__56363\,
            I => \N__56306\
        );

    \I__13958\ : InMux
    port map (
            O => \N__56362\,
            I => \N__56292\
        );

    \I__13957\ : InMux
    port map (
            O => \N__56361\,
            I => \N__56288\
        );

    \I__13956\ : InMux
    port map (
            O => \N__56360\,
            I => \N__56283\
        );

    \I__13955\ : InMux
    port map (
            O => \N__56359\,
            I => \N__56278\
        );

    \I__13954\ : InMux
    port map (
            O => \N__56358\,
            I => \N__56275\
        );

    \I__13953\ : InMux
    port map (
            O => \N__56357\,
            I => \N__56272\
        );

    \I__13952\ : LocalMux
    port map (
            O => \N__56348\,
            I => \N__56265\
        );

    \I__13951\ : LocalMux
    port map (
            O => \N__56345\,
            I => \N__56260\
        );

    \I__13950\ : LocalMux
    port map (
            O => \N__56342\,
            I => \N__56257\
        );

    \I__13949\ : InMux
    port map (
            O => \N__56341\,
            I => \N__56254\
        );

    \I__13948\ : InMux
    port map (
            O => \N__56340\,
            I => \N__56241\
        );

    \I__13947\ : InMux
    port map (
            O => \N__56339\,
            I => \N__56238\
        );

    \I__13946\ : InMux
    port map (
            O => \N__56338\,
            I => \N__56231\
        );

    \I__13945\ : InMux
    port map (
            O => \N__56337\,
            I => \N__56231\
        );

    \I__13944\ : InMux
    port map (
            O => \N__56336\,
            I => \N__56226\
        );

    \I__13943\ : InMux
    port map (
            O => \N__56335\,
            I => \N__56226\
        );

    \I__13942\ : InMux
    port map (
            O => \N__56334\,
            I => \N__56223\
        );

    \I__13941\ : InMux
    port map (
            O => \N__56333\,
            I => \N__56216\
        );

    \I__13940\ : InMux
    port map (
            O => \N__56332\,
            I => \N__56216\
        );

    \I__13939\ : InMux
    port map (
            O => \N__56331\,
            I => \N__56216\
        );

    \I__13938\ : InMux
    port map (
            O => \N__56330\,
            I => \N__56213\
        );

    \I__13937\ : InMux
    port map (
            O => \N__56329\,
            I => \N__56210\
        );

    \I__13936\ : LocalMux
    port map (
            O => \N__56326\,
            I => \N__56207\
        );

    \I__13935\ : InMux
    port map (
            O => \N__56325\,
            I => \N__56204\
        );

    \I__13934\ : InMux
    port map (
            O => \N__56324\,
            I => \N__56197\
        );

    \I__13933\ : InMux
    port map (
            O => \N__56323\,
            I => \N__56197\
        );

    \I__13932\ : InMux
    port map (
            O => \N__56322\,
            I => \N__56197\
        );

    \I__13931\ : InMux
    port map (
            O => \N__56321\,
            I => \N__56188\
        );

    \I__13930\ : InMux
    port map (
            O => \N__56320\,
            I => \N__56188\
        );

    \I__13929\ : InMux
    port map (
            O => \N__56319\,
            I => \N__56188\
        );

    \I__13928\ : InMux
    port map (
            O => \N__56318\,
            I => \N__56188\
        );

    \I__13927\ : InMux
    port map (
            O => \N__56317\,
            I => \N__56177\
        );

    \I__13926\ : LocalMux
    port map (
            O => \N__56314\,
            I => \N__56174\
        );

    \I__13925\ : InMux
    port map (
            O => \N__56313\,
            I => \N__56171\
        );

    \I__13924\ : Span4Mux_h
    port map (
            O => \N__56310\,
            I => \N__56168\
        );

    \I__13923\ : InMux
    port map (
            O => \N__56309\,
            I => \N__56163\
        );

    \I__13922\ : LocalMux
    port map (
            O => \N__56306\,
            I => \N__56160\
        );

    \I__13921\ : InMux
    port map (
            O => \N__56305\,
            I => \N__56154\
        );

    \I__13920\ : InMux
    port map (
            O => \N__56304\,
            I => \N__56154\
        );

    \I__13919\ : InMux
    port map (
            O => \N__56303\,
            I => \N__56145\
        );

    \I__13918\ : InMux
    port map (
            O => \N__56302\,
            I => \N__56145\
        );

    \I__13917\ : InMux
    port map (
            O => \N__56301\,
            I => \N__56145\
        );

    \I__13916\ : InMux
    port map (
            O => \N__56300\,
            I => \N__56145\
        );

    \I__13915\ : InMux
    port map (
            O => \N__56299\,
            I => \N__56140\
        );

    \I__13914\ : InMux
    port map (
            O => \N__56298\,
            I => \N__56137\
        );

    \I__13913\ : InMux
    port map (
            O => \N__56297\,
            I => \N__56132\
        );

    \I__13912\ : InMux
    port map (
            O => \N__56296\,
            I => \N__56132\
        );

    \I__13911\ : InMux
    port map (
            O => \N__56295\,
            I => \N__56129\
        );

    \I__13910\ : LocalMux
    port map (
            O => \N__56292\,
            I => \N__56126\
        );

    \I__13909\ : InMux
    port map (
            O => \N__56291\,
            I => \N__56123\
        );

    \I__13908\ : LocalMux
    port map (
            O => \N__56288\,
            I => \N__56120\
        );

    \I__13907\ : InMux
    port map (
            O => \N__56287\,
            I => \N__56115\
        );

    \I__13906\ : InMux
    port map (
            O => \N__56286\,
            I => \N__56115\
        );

    \I__13905\ : LocalMux
    port map (
            O => \N__56283\,
            I => \N__56112\
        );

    \I__13904\ : InMux
    port map (
            O => \N__56282\,
            I => \N__56107\
        );

    \I__13903\ : InMux
    port map (
            O => \N__56281\,
            I => \N__56107\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__56278\,
            I => \N__56103\
        );

    \I__13901\ : LocalMux
    port map (
            O => \N__56275\,
            I => \N__56100\
        );

    \I__13900\ : LocalMux
    port map (
            O => \N__56272\,
            I => \N__56097\
        );

    \I__13899\ : InMux
    port map (
            O => \N__56271\,
            I => \N__56094\
        );

    \I__13898\ : InMux
    port map (
            O => \N__56270\,
            I => \N__56087\
        );

    \I__13897\ : InMux
    port map (
            O => \N__56269\,
            I => \N__56087\
        );

    \I__13896\ : InMux
    port map (
            O => \N__56268\,
            I => \N__56087\
        );

    \I__13895\ : Span4Mux_h
    port map (
            O => \N__56265\,
            I => \N__56084\
        );

    \I__13894\ : InMux
    port map (
            O => \N__56264\,
            I => \N__56079\
        );

    \I__13893\ : InMux
    port map (
            O => \N__56263\,
            I => \N__56079\
        );

    \I__13892\ : Span4Mux_v
    port map (
            O => \N__56260\,
            I => \N__56074\
        );

    \I__13891\ : Span4Mux_h
    port map (
            O => \N__56257\,
            I => \N__56074\
        );

    \I__13890\ : LocalMux
    port map (
            O => \N__56254\,
            I => \N__56068\
        );

    \I__13889\ : InMux
    port map (
            O => \N__56253\,
            I => \N__56061\
        );

    \I__13888\ : InMux
    port map (
            O => \N__56252\,
            I => \N__56061\
        );

    \I__13887\ : InMux
    port map (
            O => \N__56251\,
            I => \N__56061\
        );

    \I__13886\ : InMux
    port map (
            O => \N__56250\,
            I => \N__56056\
        );

    \I__13885\ : InMux
    port map (
            O => \N__56249\,
            I => \N__56056\
        );

    \I__13884\ : InMux
    port map (
            O => \N__56248\,
            I => \N__56051\
        );

    \I__13883\ : InMux
    port map (
            O => \N__56247\,
            I => \N__56051\
        );

    \I__13882\ : InMux
    port map (
            O => \N__56246\,
            I => \N__56046\
        );

    \I__13881\ : InMux
    port map (
            O => \N__56245\,
            I => \N__56046\
        );

    \I__13880\ : InMux
    port map (
            O => \N__56244\,
            I => \N__56043\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__56241\,
            I => \N__56040\
        );

    \I__13878\ : LocalMux
    port map (
            O => \N__56238\,
            I => \N__56037\
        );

    \I__13877\ : InMux
    port map (
            O => \N__56237\,
            I => \N__56032\
        );

    \I__13876\ : InMux
    port map (
            O => \N__56236\,
            I => \N__56032\
        );

    \I__13875\ : LocalMux
    port map (
            O => \N__56231\,
            I => \N__56029\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__56226\,
            I => \N__56020\
        );

    \I__13873\ : LocalMux
    port map (
            O => \N__56223\,
            I => \N__56020\
        );

    \I__13872\ : LocalMux
    port map (
            O => \N__56216\,
            I => \N__56020\
        );

    \I__13871\ : LocalMux
    port map (
            O => \N__56213\,
            I => \N__56020\
        );

    \I__13870\ : LocalMux
    port map (
            O => \N__56210\,
            I => \N__56009\
        );

    \I__13869\ : Span4Mux_v
    port map (
            O => \N__56207\,
            I => \N__56009\
        );

    \I__13868\ : LocalMux
    port map (
            O => \N__56204\,
            I => \N__56009\
        );

    \I__13867\ : LocalMux
    port map (
            O => \N__56197\,
            I => \N__56009\
        );

    \I__13866\ : LocalMux
    port map (
            O => \N__56188\,
            I => \N__56009\
        );

    \I__13865\ : InMux
    port map (
            O => \N__56187\,
            I => \N__55999\
        );

    \I__13864\ : InMux
    port map (
            O => \N__56186\,
            I => \N__55999\
        );

    \I__13863\ : InMux
    port map (
            O => \N__56185\,
            I => \N__55999\
        );

    \I__13862\ : InMux
    port map (
            O => \N__56184\,
            I => \N__55996\
        );

    \I__13861\ : InMux
    port map (
            O => \N__56183\,
            I => \N__55993\
        );

    \I__13860\ : InMux
    port map (
            O => \N__56182\,
            I => \N__55988\
        );

    \I__13859\ : InMux
    port map (
            O => \N__56181\,
            I => \N__55988\
        );

    \I__13858\ : InMux
    port map (
            O => \N__56180\,
            I => \N__55985\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__56177\,
            I => \N__55978\
        );

    \I__13856\ : Span4Mux_h
    port map (
            O => \N__56174\,
            I => \N__55978\
        );

    \I__13855\ : LocalMux
    port map (
            O => \N__56171\,
            I => \N__55978\
        );

    \I__13854\ : Span4Mux_v
    port map (
            O => \N__56168\,
            I => \N__55975\
        );

    \I__13853\ : InMux
    port map (
            O => \N__56167\,
            I => \N__55970\
        );

    \I__13852\ : InMux
    port map (
            O => \N__56166\,
            I => \N__55970\
        );

    \I__13851\ : LocalMux
    port map (
            O => \N__56163\,
            I => \N__55967\
        );

    \I__13850\ : Span4Mux_h
    port map (
            O => \N__56160\,
            I => \N__55964\
        );

    \I__13849\ : InMux
    port map (
            O => \N__56159\,
            I => \N__55961\
        );

    \I__13848\ : LocalMux
    port map (
            O => \N__56154\,
            I => \N__55956\
        );

    \I__13847\ : LocalMux
    port map (
            O => \N__56145\,
            I => \N__55956\
        );

    \I__13846\ : InMux
    port map (
            O => \N__56144\,
            I => \N__55953\
        );

    \I__13845\ : InMux
    port map (
            O => \N__56143\,
            I => \N__55950\
        );

    \I__13844\ : LocalMux
    port map (
            O => \N__56140\,
            I => \N__55940\
        );

    \I__13843\ : LocalMux
    port map (
            O => \N__56137\,
            I => \N__55935\
        );

    \I__13842\ : LocalMux
    port map (
            O => \N__56132\,
            I => \N__55935\
        );

    \I__13841\ : LocalMux
    port map (
            O => \N__56129\,
            I => \N__55932\
        );

    \I__13840\ : Span4Mux_h
    port map (
            O => \N__56126\,
            I => \N__55929\
        );

    \I__13839\ : LocalMux
    port map (
            O => \N__56123\,
            I => \N__55924\
        );

    \I__13838\ : Span4Mux_h
    port map (
            O => \N__56120\,
            I => \N__55924\
        );

    \I__13837\ : LocalMux
    port map (
            O => \N__56115\,
            I => \N__55917\
        );

    \I__13836\ : Span4Mux_v
    port map (
            O => \N__56112\,
            I => \N__55917\
        );

    \I__13835\ : LocalMux
    port map (
            O => \N__56107\,
            I => \N__55917\
        );

    \I__13834\ : InMux
    port map (
            O => \N__56106\,
            I => \N__55914\
        );

    \I__13833\ : Span4Mux_h
    port map (
            O => \N__56103\,
            I => \N__55909\
        );

    \I__13832\ : Span4Mux_h
    port map (
            O => \N__56100\,
            I => \N__55909\
        );

    \I__13831\ : Span4Mux_h
    port map (
            O => \N__56097\,
            I => \N__55900\
        );

    \I__13830\ : LocalMux
    port map (
            O => \N__56094\,
            I => \N__55900\
        );

    \I__13829\ : LocalMux
    port map (
            O => \N__56087\,
            I => \N__55900\
        );

    \I__13828\ : Span4Mux_v
    port map (
            O => \N__56084\,
            I => \N__55900\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__56079\,
            I => \N__55897\
        );

    \I__13826\ : Span4Mux_v
    port map (
            O => \N__56074\,
            I => \N__55894\
        );

    \I__13825\ : InMux
    port map (
            O => \N__56073\,
            I => \N__55891\
        );

    \I__13824\ : InMux
    port map (
            O => \N__56072\,
            I => \N__55886\
        );

    \I__13823\ : InMux
    port map (
            O => \N__56071\,
            I => \N__55886\
        );

    \I__13822\ : Span4Mux_v
    port map (
            O => \N__56068\,
            I => \N__55881\
        );

    \I__13821\ : LocalMux
    port map (
            O => \N__56061\,
            I => \N__55881\
        );

    \I__13820\ : LocalMux
    port map (
            O => \N__56056\,
            I => \N__55876\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__56051\,
            I => \N__55876\
        );

    \I__13818\ : LocalMux
    port map (
            O => \N__56046\,
            I => \N__55873\
        );

    \I__13817\ : LocalMux
    port map (
            O => \N__56043\,
            I => \N__55864\
        );

    \I__13816\ : Span4Mux_h
    port map (
            O => \N__56040\,
            I => \N__55864\
        );

    \I__13815\ : Span4Mux_h
    port map (
            O => \N__56037\,
            I => \N__55864\
        );

    \I__13814\ : LocalMux
    port map (
            O => \N__56032\,
            I => \N__55864\
        );

    \I__13813\ : Span4Mux_h
    port map (
            O => \N__56029\,
            I => \N__55857\
        );

    \I__13812\ : Span4Mux_v
    port map (
            O => \N__56020\,
            I => \N__55857\
        );

    \I__13811\ : Span4Mux_v
    port map (
            O => \N__56009\,
            I => \N__55857\
        );

    \I__13810\ : InMux
    port map (
            O => \N__56008\,
            I => \N__55850\
        );

    \I__13809\ : InMux
    port map (
            O => \N__56007\,
            I => \N__55850\
        );

    \I__13808\ : InMux
    port map (
            O => \N__56006\,
            I => \N__55850\
        );

    \I__13807\ : LocalMux
    port map (
            O => \N__55999\,
            I => \N__55847\
        );

    \I__13806\ : LocalMux
    port map (
            O => \N__55996\,
            I => \N__55842\
        );

    \I__13805\ : LocalMux
    port map (
            O => \N__55993\,
            I => \N__55842\
        );

    \I__13804\ : LocalMux
    port map (
            O => \N__55988\,
            I => \N__55839\
        );

    \I__13803\ : LocalMux
    port map (
            O => \N__55985\,
            I => \N__55836\
        );

    \I__13802\ : Span4Mux_v
    port map (
            O => \N__55978\,
            I => \N__55831\
        );

    \I__13801\ : Span4Mux_v
    port map (
            O => \N__55975\,
            I => \N__55831\
        );

    \I__13800\ : LocalMux
    port map (
            O => \N__55970\,
            I => \N__55818\
        );

    \I__13799\ : Span4Mux_v
    port map (
            O => \N__55967\,
            I => \N__55818\
        );

    \I__13798\ : Span4Mux_v
    port map (
            O => \N__55964\,
            I => \N__55818\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__55961\,
            I => \N__55818\
        );

    \I__13796\ : Span4Mux_h
    port map (
            O => \N__55956\,
            I => \N__55818\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__55953\,
            I => \N__55818\
        );

    \I__13794\ : LocalMux
    port map (
            O => \N__55950\,
            I => \N__55813\
        );

    \I__13793\ : InMux
    port map (
            O => \N__55949\,
            I => \N__55810\
        );

    \I__13792\ : InMux
    port map (
            O => \N__55948\,
            I => \N__55803\
        );

    \I__13791\ : InMux
    port map (
            O => \N__55947\,
            I => \N__55803\
        );

    \I__13790\ : InMux
    port map (
            O => \N__55946\,
            I => \N__55803\
        );

    \I__13789\ : InMux
    port map (
            O => \N__55945\,
            I => \N__55798\
        );

    \I__13788\ : InMux
    port map (
            O => \N__55944\,
            I => \N__55798\
        );

    \I__13787\ : InMux
    port map (
            O => \N__55943\,
            I => \N__55795\
        );

    \I__13786\ : Span12Mux_h
    port map (
            O => \N__55940\,
            I => \N__55788\
        );

    \I__13785\ : Span12Mux_h
    port map (
            O => \N__55935\,
            I => \N__55788\
        );

    \I__13784\ : Span12Mux_h
    port map (
            O => \N__55932\,
            I => \N__55788\
        );

    \I__13783\ : Span4Mux_h
    port map (
            O => \N__55929\,
            I => \N__55781\
        );

    \I__13782\ : Span4Mux_v
    port map (
            O => \N__55924\,
            I => \N__55781\
        );

    \I__13781\ : Span4Mux_h
    port map (
            O => \N__55917\,
            I => \N__55781\
        );

    \I__13780\ : LocalMux
    port map (
            O => \N__55914\,
            I => \N__55770\
        );

    \I__13779\ : Span4Mux_v
    port map (
            O => \N__55909\,
            I => \N__55770\
        );

    \I__13778\ : Span4Mux_h
    port map (
            O => \N__55900\,
            I => \N__55770\
        );

    \I__13777\ : Span4Mux_h
    port map (
            O => \N__55897\,
            I => \N__55770\
        );

    \I__13776\ : Span4Mux_h
    port map (
            O => \N__55894\,
            I => \N__55770\
        );

    \I__13775\ : LocalMux
    port map (
            O => \N__55891\,
            I => \N__55755\
        );

    \I__13774\ : LocalMux
    port map (
            O => \N__55886\,
            I => \N__55755\
        );

    \I__13773\ : Span4Mux_v
    port map (
            O => \N__55881\,
            I => \N__55755\
        );

    \I__13772\ : Span4Mux_h
    port map (
            O => \N__55876\,
            I => \N__55755\
        );

    \I__13771\ : Span4Mux_h
    port map (
            O => \N__55873\,
            I => \N__55755\
        );

    \I__13770\ : Span4Mux_v
    port map (
            O => \N__55864\,
            I => \N__55755\
        );

    \I__13769\ : Span4Mux_h
    port map (
            O => \N__55857\,
            I => \N__55755\
        );

    \I__13768\ : LocalMux
    port map (
            O => \N__55850\,
            I => \N__55740\
        );

    \I__13767\ : Span4Mux_v
    port map (
            O => \N__55847\,
            I => \N__55740\
        );

    \I__13766\ : Span4Mux_v
    port map (
            O => \N__55842\,
            I => \N__55740\
        );

    \I__13765\ : Span4Mux_h
    port map (
            O => \N__55839\,
            I => \N__55740\
        );

    \I__13764\ : Span4Mux_h
    port map (
            O => \N__55836\,
            I => \N__55740\
        );

    \I__13763\ : Span4Mux_h
    port map (
            O => \N__55831\,
            I => \N__55740\
        );

    \I__13762\ : Span4Mux_v
    port map (
            O => \N__55818\,
            I => \N__55740\
        );

    \I__13761\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55735\
        );

    \I__13760\ : InMux
    port map (
            O => \N__55816\,
            I => \N__55735\
        );

    \I__13759\ : Odrv4
    port map (
            O => \N__55813\,
            I => comm_cmd_0
        );

    \I__13758\ : LocalMux
    port map (
            O => \N__55810\,
            I => comm_cmd_0
        );

    \I__13757\ : LocalMux
    port map (
            O => \N__55803\,
            I => comm_cmd_0
        );

    \I__13756\ : LocalMux
    port map (
            O => \N__55798\,
            I => comm_cmd_0
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__55795\,
            I => comm_cmd_0
        );

    \I__13754\ : Odrv12
    port map (
            O => \N__55788\,
            I => comm_cmd_0
        );

    \I__13753\ : Odrv4
    port map (
            O => \N__55781\,
            I => comm_cmd_0
        );

    \I__13752\ : Odrv4
    port map (
            O => \N__55770\,
            I => comm_cmd_0
        );

    \I__13751\ : Odrv4
    port map (
            O => \N__55755\,
            I => comm_cmd_0
        );

    \I__13750\ : Odrv4
    port map (
            O => \N__55740\,
            I => comm_cmd_0
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__55735\,
            I => comm_cmd_0
        );

    \I__13748\ : InMux
    port map (
            O => \N__55712\,
            I => \N__55709\
        );

    \I__13747\ : LocalMux
    port map (
            O => \N__55709\,
            I => \N__55706\
        );

    \I__13746\ : Span4Mux_h
    port map (
            O => \N__55706\,
            I => \N__55703\
        );

    \I__13745\ : Odrv4
    port map (
            O => \N__55703\,
            I => buf_data_iac_10
        );

    \I__13744\ : CascadeMux
    port map (
            O => \N__55700\,
            I => \N__55697\
        );

    \I__13743\ : InMux
    port map (
            O => \N__55697\,
            I => \N__55694\
        );

    \I__13742\ : LocalMux
    port map (
            O => \N__55694\,
            I => \N__55691\
        );

    \I__13741\ : Span4Mux_h
    port map (
            O => \N__55691\,
            I => \N__55688\
        );

    \I__13740\ : Odrv4
    port map (
            O => \N__55688\,
            I => n21320
        );

    \I__13739\ : InMux
    port map (
            O => \N__55685\,
            I => \N__55681\
        );

    \I__13738\ : InMux
    port map (
            O => \N__55684\,
            I => \N__55678\
        );

    \I__13737\ : LocalMux
    port map (
            O => \N__55681\,
            I => \N__55673\
        );

    \I__13736\ : LocalMux
    port map (
            O => \N__55678\,
            I => \N__55673\
        );

    \I__13735\ : Odrv12
    port map (
            O => \N__55673\,
            I => \comm_spi.n14655\
        );

    \I__13734\ : SRMux
    port map (
            O => \N__55670\,
            I => \N__55667\
        );

    \I__13733\ : LocalMux
    port map (
            O => \N__55667\,
            I => \N__55664\
        );

    \I__13732\ : Span4Mux_h
    port map (
            O => \N__55664\,
            I => \N__55661\
        );

    \I__13731\ : Span4Mux_v
    port map (
            O => \N__55661\,
            I => \N__55658\
        );

    \I__13730\ : Odrv4
    port map (
            O => \N__55658\,
            I => \comm_spi.data_tx_7__N_778\
        );

    \I__13729\ : InMux
    port map (
            O => \N__55655\,
            I => \N__55650\
        );

    \I__13728\ : InMux
    port map (
            O => \N__55654\,
            I => \N__55647\
        );

    \I__13727\ : InMux
    port map (
            O => \N__55653\,
            I => \N__55644\
        );

    \I__13726\ : LocalMux
    port map (
            O => \N__55650\,
            I => \comm_spi.n22673\
        );

    \I__13725\ : LocalMux
    port map (
            O => \N__55647\,
            I => \comm_spi.n22673\
        );

    \I__13724\ : LocalMux
    port map (
            O => \N__55644\,
            I => \comm_spi.n22673\
        );

    \I__13723\ : InMux
    port map (
            O => \N__55637\,
            I => \N__55633\
        );

    \I__13722\ : InMux
    port map (
            O => \N__55636\,
            I => \N__55630\
        );

    \I__13721\ : LocalMux
    port map (
            O => \N__55633\,
            I => \N__55627\
        );

    \I__13720\ : LocalMux
    port map (
            O => \N__55630\,
            I => \N__55624\
        );

    \I__13719\ : Odrv4
    port map (
            O => \N__55627\,
            I => \comm_spi.n14651\
        );

    \I__13718\ : Odrv4
    port map (
            O => \N__55624\,
            I => \comm_spi.n14651\
        );

    \I__13717\ : InMux
    port map (
            O => \N__55619\,
            I => \N__55615\
        );

    \I__13716\ : InMux
    port map (
            O => \N__55618\,
            I => \N__55612\
        );

    \I__13715\ : LocalMux
    port map (
            O => \N__55615\,
            I => \N__55607\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__55612\,
            I => \N__55607\
        );

    \I__13713\ : Odrv12
    port map (
            O => \N__55607\,
            I => \comm_spi.n14654\
        );

    \I__13712\ : SRMux
    port map (
            O => \N__55604\,
            I => \N__55601\
        );

    \I__13711\ : LocalMux
    port map (
            O => \N__55601\,
            I => \N__55598\
        );

    \I__13710\ : Span4Mux_h
    port map (
            O => \N__55598\,
            I => \N__55595\
        );

    \I__13709\ : Odrv4
    port map (
            O => \N__55595\,
            I => \comm_spi.data_tx_7__N_781\
        );

    \I__13708\ : InMux
    port map (
            O => \N__55592\,
            I => \N__55589\
        );

    \I__13707\ : LocalMux
    port map (
            O => \N__55589\,
            I => buf_data_iac_23
        );

    \I__13706\ : InMux
    port map (
            O => \N__55586\,
            I => \N__55583\
        );

    \I__13705\ : LocalMux
    port map (
            O => \N__55583\,
            I => \N__55580\
        );

    \I__13704\ : Span4Mux_v
    port map (
            O => \N__55580\,
            I => \N__55577\
        );

    \I__13703\ : Span4Mux_h
    port map (
            O => \N__55577\,
            I => \N__55574\
        );

    \I__13702\ : Span4Mux_h
    port map (
            O => \N__55574\,
            I => \N__55571\
        );

    \I__13701\ : Sp12to4
    port map (
            O => \N__55571\,
            I => \N__55568\
        );

    \I__13700\ : Odrv12
    port map (
            O => \N__55568\,
            I => n21204
        );

    \I__13699\ : IoInMux
    port map (
            O => \N__55565\,
            I => \N__55562\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__55562\,
            I => \N__55559\
        );

    \I__13697\ : Span4Mux_s3_h
    port map (
            O => \N__55559\,
            I => \N__55556\
        );

    \I__13696\ : Span4Mux_v
    port map (
            O => \N__55556\,
            I => \N__55553\
        );

    \I__13695\ : Span4Mux_v
    port map (
            O => \N__55553\,
            I => \N__55550\
        );

    \I__13694\ : Span4Mux_h
    port map (
            O => \N__55550\,
            I => \N__55547\
        );

    \I__13693\ : Odrv4
    port map (
            O => \N__55547\,
            I => \ICE_SPI_MISO\
        );

    \I__13692\ : InMux
    port map (
            O => \N__55544\,
            I => \N__55541\
        );

    \I__13691\ : LocalMux
    port map (
            O => \N__55541\,
            I => \comm_spi.n14621\
        );

    \I__13690\ : InMux
    port map (
            O => \N__55538\,
            I => \N__55535\
        );

    \I__13689\ : LocalMux
    port map (
            O => \N__55535\,
            I => \N__55531\
        );

    \I__13688\ : InMux
    port map (
            O => \N__55534\,
            I => \N__55528\
        );

    \I__13687\ : Span4Mux_h
    port map (
            O => \N__55531\,
            I => \N__55523\
        );

    \I__13686\ : LocalMux
    port map (
            O => \N__55528\,
            I => \N__55523\
        );

    \I__13685\ : Odrv4
    port map (
            O => \N__55523\,
            I => \comm_spi.n14626\
        );

    \I__13684\ : InMux
    port map (
            O => \N__55520\,
            I => \N__55517\
        );

    \I__13683\ : LocalMux
    port map (
            O => \N__55517\,
            I => \N__55514\
        );

    \I__13682\ : Odrv4
    port map (
            O => \N__55514\,
            I => \comm_spi.n14620\
        );

    \I__13681\ : InMux
    port map (
            O => \N__55511\,
            I => \N__55507\
        );

    \I__13680\ : InMux
    port map (
            O => \N__55510\,
            I => \N__55504\
        );

    \I__13679\ : LocalMux
    port map (
            O => \N__55507\,
            I => \N__55501\
        );

    \I__13678\ : LocalMux
    port map (
            O => \N__55504\,
            I => \N__55498\
        );

    \I__13677\ : Span4Mux_v
    port map (
            O => \N__55501\,
            I => \N__55492\
        );

    \I__13676\ : Span4Mux_h
    port map (
            O => \N__55498\,
            I => \N__55492\
        );

    \I__13675\ : InMux
    port map (
            O => \N__55497\,
            I => \N__55489\
        );

    \I__13674\ : Span4Mux_v
    port map (
            O => \N__55492\,
            I => \N__55484\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__55489\,
            I => \N__55484\
        );

    \I__13672\ : Span4Mux_v
    port map (
            O => \N__55484\,
            I => \N__55481\
        );

    \I__13671\ : Odrv4
    port map (
            O => \N__55481\,
            I => comm_tx_buf_6
        );

    \I__13670\ : InMux
    port map (
            O => \N__55478\,
            I => \N__55473\
        );

    \I__13669\ : InMux
    port map (
            O => \N__55477\,
            I => \N__55470\
        );

    \I__13668\ : InMux
    port map (
            O => \N__55476\,
            I => \N__55466\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__55473\,
            I => \N__55460\
        );

    \I__13666\ : LocalMux
    port map (
            O => \N__55470\,
            I => \N__55460\
        );

    \I__13665\ : InMux
    port map (
            O => \N__55469\,
            I => \N__55457\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__55466\,
            I => \N__55454\
        );

    \I__13663\ : InMux
    port map (
            O => \N__55465\,
            I => \N__55451\
        );

    \I__13662\ : Span4Mux_v
    port map (
            O => \N__55460\,
            I => \N__55445\
        );

    \I__13661\ : LocalMux
    port map (
            O => \N__55457\,
            I => \N__55445\
        );

    \I__13660\ : Span4Mux_v
    port map (
            O => \N__55454\,
            I => \N__55440\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__55451\,
            I => \N__55440\
        );

    \I__13658\ : InMux
    port map (
            O => \N__55450\,
            I => \N__55437\
        );

    \I__13657\ : Span4Mux_h
    port map (
            O => \N__55445\,
            I => \N__55434\
        );

    \I__13656\ : Odrv4
    port map (
            O => \N__55440\,
            I => \comm_spi.n14619\
        );

    \I__13655\ : LocalMux
    port map (
            O => \N__55437\,
            I => \comm_spi.n14619\
        );

    \I__13654\ : Odrv4
    port map (
            O => \N__55434\,
            I => \comm_spi.n14619\
        );

    \I__13653\ : InMux
    port map (
            O => \N__55427\,
            I => \N__55424\
        );

    \I__13652\ : LocalMux
    port map (
            O => \N__55424\,
            I => \N__55420\
        );

    \I__13651\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55417\
        );

    \I__13650\ : Odrv4
    port map (
            O => \N__55420\,
            I => \comm_spi.n14627\
        );

    \I__13649\ : LocalMux
    port map (
            O => \N__55417\,
            I => \comm_spi.n14627\
        );

    \I__13648\ : InMux
    port map (
            O => \N__55412\,
            I => \N__55408\
        );

    \I__13647\ : InMux
    port map (
            O => \N__55411\,
            I => \N__55405\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__55408\,
            I => \comm_spi.n14624\
        );

    \I__13645\ : LocalMux
    port map (
            O => \N__55405\,
            I => \comm_spi.n14624\
        );

    \I__13644\ : InMux
    port map (
            O => \N__55400\,
            I => \N__55397\
        );

    \I__13643\ : LocalMux
    port map (
            O => \N__55397\,
            I => \N__55394\
        );

    \I__13642\ : Span4Mux_v
    port map (
            O => \N__55394\,
            I => \N__55390\
        );

    \I__13641\ : InMux
    port map (
            O => \N__55393\,
            I => \N__55387\
        );

    \I__13640\ : Span4Mux_h
    port map (
            O => \N__55390\,
            I => \N__55381\
        );

    \I__13639\ : LocalMux
    port map (
            O => \N__55387\,
            I => \N__55381\
        );

    \I__13638\ : InMux
    port map (
            O => \N__55386\,
            I => \N__55378\
        );

    \I__13637\ : Odrv4
    port map (
            O => \N__55381\,
            I => \comm_spi.n22682\
        );

    \I__13636\ : LocalMux
    port map (
            O => \N__55378\,
            I => \comm_spi.n22682\
        );

    \I__13635\ : InMux
    port map (
            O => \N__55373\,
            I => \N__55370\
        );

    \I__13634\ : LocalMux
    port map (
            O => \N__55370\,
            I => \N__55367\
        );

    \I__13633\ : Sp12to4
    port map (
            O => \N__55367\,
            I => \N__55363\
        );

    \I__13632\ : InMux
    port map (
            O => \N__55366\,
            I => \N__55360\
        );

    \I__13631\ : Span12Mux_h
    port map (
            O => \N__55363\,
            I => \N__55357\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__55360\,
            I => \N__55354\
        );

    \I__13629\ : Odrv12
    port map (
            O => \N__55357\,
            I => \comm_spi.n14638\
        );

    \I__13628\ : Odrv4
    port map (
            O => \N__55354\,
            I => \comm_spi.n14638\
        );

    \I__13627\ : InMux
    port map (
            O => \N__55349\,
            I => \N__55346\
        );

    \I__13626\ : LocalMux
    port map (
            O => \N__55346\,
            I => \N__55343\
        );

    \I__13625\ : Span4Mux_h
    port map (
            O => \N__55343\,
            I => \N__55340\
        );

    \I__13624\ : Span4Mux_h
    port map (
            O => \N__55340\,
            I => \N__55336\
        );

    \I__13623\ : InMux
    port map (
            O => \N__55339\,
            I => \N__55333\
        );

    \I__13622\ : Sp12to4
    port map (
            O => \N__55336\,
            I => \N__55328\
        );

    \I__13621\ : LocalMux
    port map (
            O => \N__55333\,
            I => \N__55328\
        );

    \I__13620\ : Odrv12
    port map (
            O => \N__55328\,
            I => \comm_spi.n14639\
        );

    \I__13619\ : SRMux
    port map (
            O => \N__55325\,
            I => \N__55322\
        );

    \I__13618\ : LocalMux
    port map (
            O => \N__55322\,
            I => \comm_spi.data_tx_7__N_787\
        );

    \I__13617\ : InMux
    port map (
            O => \N__55319\,
            I => \N__55315\
        );

    \I__13616\ : InMux
    port map (
            O => \N__55318\,
            I => \N__55312\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__55315\,
            I => \N__55308\
        );

    \I__13614\ : LocalMux
    port map (
            O => \N__55312\,
            I => \N__55305\
        );

    \I__13613\ : InMux
    port map (
            O => \N__55311\,
            I => \N__55302\
        );

    \I__13612\ : Span4Mux_v
    port map (
            O => \N__55308\,
            I => \N__55299\
        );

    \I__13611\ : Span4Mux_v
    port map (
            O => \N__55305\,
            I => \N__55294\
        );

    \I__13610\ : LocalMux
    port map (
            O => \N__55302\,
            I => \N__55294\
        );

    \I__13609\ : Sp12to4
    port map (
            O => \N__55299\,
            I => \N__55291\
        );

    \I__13608\ : Span4Mux_h
    port map (
            O => \N__55294\,
            I => \N__55288\
        );

    \I__13607\ : Span12Mux_h
    port map (
            O => \N__55291\,
            I => \N__55283\
        );

    \I__13606\ : Sp12to4
    port map (
            O => \N__55288\,
            I => \N__55283\
        );

    \I__13605\ : Odrv12
    port map (
            O => \N__55283\,
            I => comm_tx_buf_3
        );

    \I__13604\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55276\
        );

    \I__13603\ : InMux
    port map (
            O => \N__55279\,
            I => \N__55273\
        );

    \I__13602\ : LocalMux
    port map (
            O => \N__55276\,
            I => \N__55267\
        );

    \I__13601\ : LocalMux
    port map (
            O => \N__55273\,
            I => \N__55267\
        );

    \I__13600\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55264\
        );

    \I__13599\ : Span4Mux_v
    port map (
            O => \N__55267\,
            I => \N__55259\
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__55264\,
            I => \N__55259\
        );

    \I__13597\ : Span4Mux_v
    port map (
            O => \N__55259\,
            I => \N__55256\
        );

    \I__13596\ : Span4Mux_v
    port map (
            O => \N__55256\,
            I => \N__55253\
        );

    \I__13595\ : Span4Mux_h
    port map (
            O => \N__55253\,
            I => \N__55250\
        );

    \I__13594\ : Odrv4
    port map (
            O => \N__55250\,
            I => comm_tx_buf_4
        );

    \I__13593\ : InMux
    port map (
            O => \N__55247\,
            I => \N__55241\
        );

    \I__13592\ : InMux
    port map (
            O => \N__55246\,
            I => \N__55241\
        );

    \I__13591\ : LocalMux
    port map (
            O => \N__55241\,
            I => \N__55238\
        );

    \I__13590\ : Span4Mux_h
    port map (
            O => \N__55238\,
            I => \N__55234\
        );

    \I__13589\ : InMux
    port map (
            O => \N__55237\,
            I => \N__55231\
        );

    \I__13588\ : Sp12to4
    port map (
            O => \N__55234\,
            I => \N__55226\
        );

    \I__13587\ : LocalMux
    port map (
            O => \N__55231\,
            I => \N__55226\
        );

    \I__13586\ : Span12Mux_v
    port map (
            O => \N__55226\,
            I => \N__55223\
        );

    \I__13585\ : Odrv12
    port map (
            O => \N__55223\,
            I => comm_tx_buf_5
        );

    \I__13584\ : InMux
    port map (
            O => \N__55220\,
            I => \N__55215\
        );

    \I__13583\ : InMux
    port map (
            O => \N__55219\,
            I => \N__55212\
        );

    \I__13582\ : InMux
    port map (
            O => \N__55218\,
            I => \N__55209\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__55215\,
            I => \comm_spi.n22679\
        );

    \I__13580\ : LocalMux
    port map (
            O => \N__55212\,
            I => \comm_spi.n22679\
        );

    \I__13579\ : LocalMux
    port map (
            O => \N__55209\,
            I => \comm_spi.n22679\
        );

    \I__13578\ : InMux
    port map (
            O => \N__55202\,
            I => \N__55198\
        );

    \I__13577\ : InMux
    port map (
            O => \N__55201\,
            I => \N__55195\
        );

    \I__13576\ : LocalMux
    port map (
            O => \N__55198\,
            I => \N__55190\
        );

    \I__13575\ : LocalMux
    port map (
            O => \N__55195\,
            I => \N__55190\
        );

    \I__13574\ : Odrv12
    port map (
            O => \N__55190\,
            I => \comm_spi.n14642\
        );

    \I__13573\ : InMux
    port map (
            O => \N__55187\,
            I => \N__55183\
        );

    \I__13572\ : InMux
    port map (
            O => \N__55186\,
            I => \N__55180\
        );

    \I__13571\ : LocalMux
    port map (
            O => \N__55183\,
            I => \N__55175\
        );

    \I__13570\ : LocalMux
    port map (
            O => \N__55180\,
            I => \N__55175\
        );

    \I__13569\ : Odrv4
    port map (
            O => \N__55175\,
            I => \comm_spi.n14643\
        );

    \I__13568\ : SRMux
    port map (
            O => \N__55172\,
            I => \N__55169\
        );

    \I__13567\ : LocalMux
    port map (
            O => \N__55169\,
            I => \N__55166\
        );

    \I__13566\ : Span4Mux_v
    port map (
            O => \N__55166\,
            I => \N__55163\
        );

    \I__13565\ : Odrv4
    port map (
            O => \N__55163\,
            I => \comm_spi.data_tx_7__N_784\
        );

    \I__13564\ : InMux
    port map (
            O => \N__55160\,
            I => \N__55157\
        );

    \I__13563\ : LocalMux
    port map (
            O => \N__55157\,
            I => \N__55154\
        );

    \I__13562\ : Span4Mux_v
    port map (
            O => \N__55154\,
            I => \N__55149\
        );

    \I__13561\ : InMux
    port map (
            O => \N__55153\,
            I => \N__55144\
        );

    \I__13560\ : InMux
    port map (
            O => \N__55152\,
            I => \N__55144\
        );

    \I__13559\ : Span4Mux_v
    port map (
            O => \N__55149\,
            I => \N__55141\
        );

    \I__13558\ : LocalMux
    port map (
            O => \N__55144\,
            I => \N__55138\
        );

    \I__13557\ : Sp12to4
    port map (
            O => \N__55141\,
            I => \N__55135\
        );

    \I__13556\ : Span4Mux_h
    port map (
            O => \N__55138\,
            I => \N__55132\
        );

    \I__13555\ : Odrv12
    port map (
            O => \N__55135\,
            I => comm_tx_buf_2
        );

    \I__13554\ : Odrv4
    port map (
            O => \N__55132\,
            I => comm_tx_buf_2
        );

    \I__13553\ : InMux
    port map (
            O => \N__55127\,
            I => \N__55124\
        );

    \I__13552\ : LocalMux
    port map (
            O => \N__55124\,
            I => \N__55120\
        );

    \I__13551\ : InMux
    port map (
            O => \N__55123\,
            I => \N__55117\
        );

    \I__13550\ : Span4Mux_v
    port map (
            O => \N__55120\,
            I => \N__55112\
        );

    \I__13549\ : LocalMux
    port map (
            O => \N__55117\,
            I => \N__55112\
        );

    \I__13548\ : Span4Mux_v
    port map (
            O => \N__55112\,
            I => \N__55109\
        );

    \I__13547\ : Odrv4
    port map (
            O => \N__55109\,
            I => \comm_spi.imosi\
        );

    \I__13546\ : SRMux
    port map (
            O => \N__55106\,
            I => \N__55103\
        );

    \I__13545\ : LocalMux
    port map (
            O => \N__55103\,
            I => \N__55100\
        );

    \I__13544\ : Span4Mux_v
    port map (
            O => \N__55100\,
            I => \N__55097\
        );

    \I__13543\ : Odrv4
    port map (
            O => \N__55097\,
            I => \comm_spi.DOUT_7__N_748\
        );

    \I__13542\ : SRMux
    port map (
            O => \N__55094\,
            I => \N__55091\
        );

    \I__13541\ : LocalMux
    port map (
            O => \N__55091\,
            I => \N__55088\
        );

    \I__13540\ : Span4Mux_h
    port map (
            O => \N__55088\,
            I => \N__55085\
        );

    \I__13539\ : Odrv4
    port map (
            O => \N__55085\,
            I => \comm_spi.imosi_N_753\
        );

    \I__13538\ : SRMux
    port map (
            O => \N__55082\,
            I => \N__55079\
        );

    \I__13537\ : LocalMux
    port map (
            O => \N__55079\,
            I => \N__55076\
        );

    \I__13536\ : Span4Mux_v
    port map (
            O => \N__55076\,
            I => \N__55073\
        );

    \I__13535\ : Odrv4
    port map (
            O => \N__55073\,
            I => \comm_spi.data_tx_7__N_790\
        );

    \I__13534\ : InMux
    port map (
            O => \N__55070\,
            I => \N__55065\
        );

    \I__13533\ : InMux
    port map (
            O => \N__55069\,
            I => \N__55062\
        );

    \I__13532\ : InMux
    port map (
            O => \N__55068\,
            I => \N__55059\
        );

    \I__13531\ : LocalMux
    port map (
            O => \N__55065\,
            I => \comm_spi.n22685\
        );

    \I__13530\ : LocalMux
    port map (
            O => \N__55062\,
            I => \comm_spi.n22685\
        );

    \I__13529\ : LocalMux
    port map (
            O => \N__55059\,
            I => \comm_spi.n22685\
        );

    \I__13528\ : SRMux
    port map (
            O => \N__55052\,
            I => \N__55049\
        );

    \I__13527\ : LocalMux
    port map (
            O => \N__55049\,
            I => \N__55046\
        );

    \I__13526\ : Odrv4
    port map (
            O => \N__55046\,
            I => \comm_spi.data_tx_7__N_772\
        );

    \I__13525\ : InMux
    port map (
            O => \N__55043\,
            I => \N__55040\
        );

    \I__13524\ : LocalMux
    port map (
            O => \N__55040\,
            I => \N__55036\
        );

    \I__13523\ : InMux
    port map (
            O => \N__55039\,
            I => \N__55033\
        );

    \I__13522\ : Odrv4
    port map (
            O => \N__55036\,
            I => \comm_spi.n14634\
        );

    \I__13521\ : LocalMux
    port map (
            O => \N__55033\,
            I => \comm_spi.n14634\
        );

    \I__13520\ : InMux
    port map (
            O => \N__55028\,
            I => \N__55024\
        );

    \I__13519\ : InMux
    port map (
            O => \N__55027\,
            I => \N__55021\
        );

    \I__13518\ : LocalMux
    port map (
            O => \N__55024\,
            I => \N__55017\
        );

    \I__13517\ : LocalMux
    port map (
            O => \N__55021\,
            I => \N__55014\
        );

    \I__13516\ : InMux
    port map (
            O => \N__55020\,
            I => \N__55011\
        );

    \I__13515\ : Span4Mux_v
    port map (
            O => \N__55017\,
            I => \N__55008\
        );

    \I__13514\ : Span4Mux_v
    port map (
            O => \N__55014\,
            I => \N__55003\
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__55011\,
            I => \N__55003\
        );

    \I__13512\ : Span4Mux_v
    port map (
            O => \N__55008\,
            I => \N__55000\
        );

    \I__13511\ : Span4Mux_v
    port map (
            O => \N__55003\,
            I => \N__54997\
        );

    \I__13510\ : Odrv4
    port map (
            O => \N__55000\,
            I => comm_tx_buf_1
        );

    \I__13509\ : Odrv4
    port map (
            O => \N__54997\,
            I => comm_tx_buf_1
        );

    \I__13508\ : SRMux
    port map (
            O => \N__54992\,
            I => \N__54989\
        );

    \I__13507\ : LocalMux
    port map (
            O => \N__54989\,
            I => \N__54986\
        );

    \I__13506\ : Odrv4
    port map (
            O => \N__54986\,
            I => \comm_spi.data_tx_7__N_773\
        );

    \I__13505\ : CascadeMux
    port map (
            O => \N__54983\,
            I => \N__54978\
        );

    \I__13504\ : InMux
    port map (
            O => \N__54982\,
            I => \N__54968\
        );

    \I__13503\ : InMux
    port map (
            O => \N__54981\,
            I => \N__54955\
        );

    \I__13502\ : InMux
    port map (
            O => \N__54978\,
            I => \N__54955\
        );

    \I__13501\ : CascadeMux
    port map (
            O => \N__54977\,
            I => \N__54950\
        );

    \I__13500\ : InMux
    port map (
            O => \N__54976\,
            I => \N__54932\
        );

    \I__13499\ : InMux
    port map (
            O => \N__54975\,
            I => \N__54932\
        );

    \I__13498\ : InMux
    port map (
            O => \N__54974\,
            I => \N__54932\
        );

    \I__13497\ : InMux
    port map (
            O => \N__54973\,
            I => \N__54932\
        );

    \I__13496\ : InMux
    port map (
            O => \N__54972\,
            I => \N__54932\
        );

    \I__13495\ : InMux
    port map (
            O => \N__54971\,
            I => \N__54932\
        );

    \I__13494\ : LocalMux
    port map (
            O => \N__54968\,
            I => \N__54929\
        );

    \I__13493\ : InMux
    port map (
            O => \N__54967\,
            I => \N__54924\
        );

    \I__13492\ : InMux
    port map (
            O => \N__54966\,
            I => \N__54924\
        );

    \I__13491\ : InMux
    port map (
            O => \N__54965\,
            I => \N__54917\
        );

    \I__13490\ : InMux
    port map (
            O => \N__54964\,
            I => \N__54917\
        );

    \I__13489\ : InMux
    port map (
            O => \N__54963\,
            I => \N__54914\
        );

    \I__13488\ : CascadeMux
    port map (
            O => \N__54962\,
            I => \N__54908\
        );

    \I__13487\ : CascadeMux
    port map (
            O => \N__54961\,
            I => \N__54904\
        );

    \I__13486\ : CascadeMux
    port map (
            O => \N__54960\,
            I => \N__54896\
        );

    \I__13485\ : LocalMux
    port map (
            O => \N__54955\,
            I => \N__54884\
        );

    \I__13484\ : InMux
    port map (
            O => \N__54954\,
            I => \N__54879\
        );

    \I__13483\ : InMux
    port map (
            O => \N__54953\,
            I => \N__54879\
        );

    \I__13482\ : InMux
    port map (
            O => \N__54950\,
            I => \N__54872\
        );

    \I__13481\ : InMux
    port map (
            O => \N__54949\,
            I => \N__54872\
        );

    \I__13480\ : InMux
    port map (
            O => \N__54948\,
            I => \N__54872\
        );

    \I__13479\ : InMux
    port map (
            O => \N__54947\,
            I => \N__54864\
        );

    \I__13478\ : InMux
    port map (
            O => \N__54946\,
            I => \N__54859\
        );

    \I__13477\ : InMux
    port map (
            O => \N__54945\,
            I => \N__54859\
        );

    \I__13476\ : LocalMux
    port map (
            O => \N__54932\,
            I => \N__54854\
        );

    \I__13475\ : Span4Mux_v
    port map (
            O => \N__54929\,
            I => \N__54854\
        );

    \I__13474\ : LocalMux
    port map (
            O => \N__54924\,
            I => \N__54851\
        );

    \I__13473\ : InMux
    port map (
            O => \N__54923\,
            I => \N__54848\
        );

    \I__13472\ : InMux
    port map (
            O => \N__54922\,
            I => \N__54843\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__54917\,
            I => \N__54838\
        );

    \I__13470\ : LocalMux
    port map (
            O => \N__54914\,
            I => \N__54838\
        );

    \I__13469\ : InMux
    port map (
            O => \N__54913\,
            I => \N__54833\
        );

    \I__13468\ : InMux
    port map (
            O => \N__54912\,
            I => \N__54830\
        );

    \I__13467\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54825\
        );

    \I__13466\ : InMux
    port map (
            O => \N__54908\,
            I => \N__54818\
        );

    \I__13465\ : InMux
    port map (
            O => \N__54907\,
            I => \N__54818\
        );

    \I__13464\ : InMux
    port map (
            O => \N__54904\,
            I => \N__54811\
        );

    \I__13463\ : InMux
    port map (
            O => \N__54903\,
            I => \N__54811\
        );

    \I__13462\ : InMux
    port map (
            O => \N__54902\,
            I => \N__54811\
        );

    \I__13461\ : InMux
    port map (
            O => \N__54901\,
            I => \N__54796\
        );

    \I__13460\ : InMux
    port map (
            O => \N__54900\,
            I => \N__54796\
        );

    \I__13459\ : InMux
    port map (
            O => \N__54899\,
            I => \N__54796\
        );

    \I__13458\ : InMux
    port map (
            O => \N__54896\,
            I => \N__54785\
        );

    \I__13457\ : InMux
    port map (
            O => \N__54895\,
            I => \N__54785\
        );

    \I__13456\ : InMux
    port map (
            O => \N__54894\,
            I => \N__54785\
        );

    \I__13455\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54785\
        );

    \I__13454\ : InMux
    port map (
            O => \N__54892\,
            I => \N__54785\
        );

    \I__13453\ : InMux
    port map (
            O => \N__54891\,
            I => \N__54776\
        );

    \I__13452\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54776\
        );

    \I__13451\ : InMux
    port map (
            O => \N__54889\,
            I => \N__54776\
        );

    \I__13450\ : InMux
    port map (
            O => \N__54888\,
            I => \N__54776\
        );

    \I__13449\ : InMux
    port map (
            O => \N__54887\,
            I => \N__54773\
        );

    \I__13448\ : Span4Mux_v
    port map (
            O => \N__54884\,
            I => \N__54766\
        );

    \I__13447\ : LocalMux
    port map (
            O => \N__54879\,
            I => \N__54766\
        );

    \I__13446\ : LocalMux
    port map (
            O => \N__54872\,
            I => \N__54766\
        );

    \I__13445\ : InMux
    port map (
            O => \N__54871\,
            I => \N__54758\
        );

    \I__13444\ : InMux
    port map (
            O => \N__54870\,
            I => \N__54758\
        );

    \I__13443\ : InMux
    port map (
            O => \N__54869\,
            I => \N__54751\
        );

    \I__13442\ : InMux
    port map (
            O => \N__54868\,
            I => \N__54751\
        );

    \I__13441\ : InMux
    port map (
            O => \N__54867\,
            I => \N__54751\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__54864\,
            I => \N__54740\
        );

    \I__13439\ : LocalMux
    port map (
            O => \N__54859\,
            I => \N__54740\
        );

    \I__13438\ : Span4Mux_v
    port map (
            O => \N__54854\,
            I => \N__54740\
        );

    \I__13437\ : Span4Mux_h
    port map (
            O => \N__54851\,
            I => \N__54740\
        );

    \I__13436\ : LocalMux
    port map (
            O => \N__54848\,
            I => \N__54740\
        );

    \I__13435\ : InMux
    port map (
            O => \N__54847\,
            I => \N__54737\
        );

    \I__13434\ : InMux
    port map (
            O => \N__54846\,
            I => \N__54732\
        );

    \I__13433\ : LocalMux
    port map (
            O => \N__54843\,
            I => \N__54727\
        );

    \I__13432\ : Span4Mux_v
    port map (
            O => \N__54838\,
            I => \N__54727\
        );

    \I__13431\ : CascadeMux
    port map (
            O => \N__54837\,
            I => \N__54724\
        );

    \I__13430\ : SRMux
    port map (
            O => \N__54836\,
            I => \N__54719\
        );

    \I__13429\ : LocalMux
    port map (
            O => \N__54833\,
            I => \N__54714\
        );

    \I__13428\ : LocalMux
    port map (
            O => \N__54830\,
            I => \N__54711\
        );

    \I__13427\ : InMux
    port map (
            O => \N__54829\,
            I => \N__54700\
        );

    \I__13426\ : InMux
    port map (
            O => \N__54828\,
            I => \N__54700\
        );

    \I__13425\ : LocalMux
    port map (
            O => \N__54825\,
            I => \N__54697\
        );

    \I__13424\ : InMux
    port map (
            O => \N__54824\,
            I => \N__54694\
        );

    \I__13423\ : InMux
    port map (
            O => \N__54823\,
            I => \N__54691\
        );

    \I__13422\ : LocalMux
    port map (
            O => \N__54818\,
            I => \N__54686\
        );

    \I__13421\ : LocalMux
    port map (
            O => \N__54811\,
            I => \N__54686\
        );

    \I__13420\ : InMux
    port map (
            O => \N__54810\,
            I => \N__54677\
        );

    \I__13419\ : InMux
    port map (
            O => \N__54809\,
            I => \N__54677\
        );

    \I__13418\ : InMux
    port map (
            O => \N__54808\,
            I => \N__54677\
        );

    \I__13417\ : InMux
    port map (
            O => \N__54807\,
            I => \N__54677\
        );

    \I__13416\ : InMux
    port map (
            O => \N__54806\,
            I => \N__54668\
        );

    \I__13415\ : InMux
    port map (
            O => \N__54805\,
            I => \N__54668\
        );

    \I__13414\ : InMux
    port map (
            O => \N__54804\,
            I => \N__54668\
        );

    \I__13413\ : InMux
    port map (
            O => \N__54803\,
            I => \N__54668\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__54796\,
            I => \N__54661\
        );

    \I__13411\ : LocalMux
    port map (
            O => \N__54785\,
            I => \N__54661\
        );

    \I__13410\ : LocalMux
    port map (
            O => \N__54776\,
            I => \N__54661\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__54773\,
            I => \N__54656\
        );

    \I__13408\ : Span4Mux_h
    port map (
            O => \N__54766\,
            I => \N__54656\
        );

    \I__13407\ : InMux
    port map (
            O => \N__54765\,
            I => \N__54649\
        );

    \I__13406\ : InMux
    port map (
            O => \N__54764\,
            I => \N__54649\
        );

    \I__13405\ : InMux
    port map (
            O => \N__54763\,
            I => \N__54646\
        );

    \I__13404\ : LocalMux
    port map (
            O => \N__54758\,
            I => \N__54641\
        );

    \I__13403\ : LocalMux
    port map (
            O => \N__54751\,
            I => \N__54641\
        );

    \I__13402\ : Span4Mux_v
    port map (
            O => \N__54740\,
            I => \N__54638\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__54737\,
            I => \N__54632\
        );

    \I__13400\ : InMux
    port map (
            O => \N__54736\,
            I => \N__54629\
        );

    \I__13399\ : InMux
    port map (
            O => \N__54735\,
            I => \N__54626\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__54732\,
            I => \N__54621\
        );

    \I__13397\ : Span4Mux_v
    port map (
            O => \N__54727\,
            I => \N__54621\
        );

    \I__13396\ : InMux
    port map (
            O => \N__54724\,
            I => \N__54616\
        );

    \I__13395\ : InMux
    port map (
            O => \N__54723\,
            I => \N__54616\
        );

    \I__13394\ : InMux
    port map (
            O => \N__54722\,
            I => \N__54613\
        );

    \I__13393\ : LocalMux
    port map (
            O => \N__54719\,
            I => \N__54610\
        );

    \I__13392\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54605\
        );

    \I__13391\ : InMux
    port map (
            O => \N__54717\,
            I => \N__54605\
        );

    \I__13390\ : Span4Mux_v
    port map (
            O => \N__54714\,
            I => \N__54600\
        );

    \I__13389\ : Span4Mux_v
    port map (
            O => \N__54711\,
            I => \N__54600\
        );

    \I__13388\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54593\
        );

    \I__13387\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54593\
        );

    \I__13386\ : InMux
    port map (
            O => \N__54708\,
            I => \N__54593\
        );

    \I__13385\ : InMux
    port map (
            O => \N__54707\,
            I => \N__54588\
        );

    \I__13384\ : InMux
    port map (
            O => \N__54706\,
            I => \N__54588\
        );

    \I__13383\ : InMux
    port map (
            O => \N__54705\,
            I => \N__54585\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__54700\,
            I => \N__54580\
        );

    \I__13381\ : Span4Mux_v
    port map (
            O => \N__54697\,
            I => \N__54580\
        );

    \I__13380\ : LocalMux
    port map (
            O => \N__54694\,
            I => \N__54577\
        );

    \I__13379\ : LocalMux
    port map (
            O => \N__54691\,
            I => \N__54566\
        );

    \I__13378\ : Span4Mux_v
    port map (
            O => \N__54686\,
            I => \N__54566\
        );

    \I__13377\ : LocalMux
    port map (
            O => \N__54677\,
            I => \N__54566\
        );

    \I__13376\ : LocalMux
    port map (
            O => \N__54668\,
            I => \N__54566\
        );

    \I__13375\ : Span4Mux_v
    port map (
            O => \N__54661\,
            I => \N__54566\
        );

    \I__13374\ : Span4Mux_h
    port map (
            O => \N__54656\,
            I => \N__54563\
        );

    \I__13373\ : InMux
    port map (
            O => \N__54655\,
            I => \N__54560\
        );

    \I__13372\ : InMux
    port map (
            O => \N__54654\,
            I => \N__54555\
        );

    \I__13371\ : LocalMux
    port map (
            O => \N__54649\,
            I => \N__54548\
        );

    \I__13370\ : LocalMux
    port map (
            O => \N__54646\,
            I => \N__54548\
        );

    \I__13369\ : Span4Mux_v
    port map (
            O => \N__54641\,
            I => \N__54548\
        );

    \I__13368\ : Span4Mux_h
    port map (
            O => \N__54638\,
            I => \N__54545\
        );

    \I__13367\ : InMux
    port map (
            O => \N__54637\,
            I => \N__54538\
        );

    \I__13366\ : InMux
    port map (
            O => \N__54636\,
            I => \N__54538\
        );

    \I__13365\ : InMux
    port map (
            O => \N__54635\,
            I => \N__54538\
        );

    \I__13364\ : Span4Mux_h
    port map (
            O => \N__54632\,
            I => \N__54534\
        );

    \I__13363\ : LocalMux
    port map (
            O => \N__54629\,
            I => \N__54531\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__54626\,
            I => \N__54525\
        );

    \I__13361\ : Span4Mux_v
    port map (
            O => \N__54621\,
            I => \N__54522\
        );

    \I__13360\ : LocalMux
    port map (
            O => \N__54616\,
            I => \N__54507\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__54613\,
            I => \N__54507\
        );

    \I__13358\ : Span4Mux_v
    port map (
            O => \N__54610\,
            I => \N__54507\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__54605\,
            I => \N__54507\
        );

    \I__13356\ : Span4Mux_v
    port map (
            O => \N__54600\,
            I => \N__54507\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__54593\,
            I => \N__54507\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__54588\,
            I => \N__54507\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__54585\,
            I => \N__54496\
        );

    \I__13352\ : Span4Mux_h
    port map (
            O => \N__54580\,
            I => \N__54496\
        );

    \I__13351\ : Span4Mux_h
    port map (
            O => \N__54577\,
            I => \N__54496\
        );

    \I__13350\ : Span4Mux_h
    port map (
            O => \N__54566\,
            I => \N__54496\
        );

    \I__13349\ : Span4Mux_v
    port map (
            O => \N__54563\,
            I => \N__54496\
        );

    \I__13348\ : LocalMux
    port map (
            O => \N__54560\,
            I => \N__54493\
        );

    \I__13347\ : InMux
    port map (
            O => \N__54559\,
            I => \N__54488\
        );

    \I__13346\ : InMux
    port map (
            O => \N__54558\,
            I => \N__54488\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__54555\,
            I => \N__54479\
        );

    \I__13344\ : Span4Mux_v
    port map (
            O => \N__54548\,
            I => \N__54479\
        );

    \I__13343\ : Span4Mux_h
    port map (
            O => \N__54545\,
            I => \N__54479\
        );

    \I__13342\ : LocalMux
    port map (
            O => \N__54538\,
            I => \N__54479\
        );

    \I__13341\ : InMux
    port map (
            O => \N__54537\,
            I => \N__54476\
        );

    \I__13340\ : Sp12to4
    port map (
            O => \N__54534\,
            I => \N__54471\
        );

    \I__13339\ : Span12Mux_s11_v
    port map (
            O => \N__54531\,
            I => \N__54471\
        );

    \I__13338\ : InMux
    port map (
            O => \N__54530\,
            I => \N__54468\
        );

    \I__13337\ : InMux
    port map (
            O => \N__54529\,
            I => \N__54463\
        );

    \I__13336\ : InMux
    port map (
            O => \N__54528\,
            I => \N__54463\
        );

    \I__13335\ : Span4Mux_v
    port map (
            O => \N__54525\,
            I => \N__54456\
        );

    \I__13334\ : Span4Mux_h
    port map (
            O => \N__54522\,
            I => \N__54456\
        );

    \I__13333\ : Span4Mux_v
    port map (
            O => \N__54507\,
            I => \N__54456\
        );

    \I__13332\ : Span4Mux_v
    port map (
            O => \N__54496\,
            I => \N__54453\
        );

    \I__13331\ : Span4Mux_v
    port map (
            O => \N__54493\,
            I => \N__54446\
        );

    \I__13330\ : LocalMux
    port map (
            O => \N__54488\,
            I => \N__54446\
        );

    \I__13329\ : Span4Mux_v
    port map (
            O => \N__54479\,
            I => \N__54446\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__54476\,
            I => comm_state_3
        );

    \I__13327\ : Odrv12
    port map (
            O => \N__54471\,
            I => comm_state_3
        );

    \I__13326\ : LocalMux
    port map (
            O => \N__54468\,
            I => comm_state_3
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__54463\,
            I => comm_state_3
        );

    \I__13324\ : Odrv4
    port map (
            O => \N__54456\,
            I => comm_state_3
        );

    \I__13323\ : Odrv4
    port map (
            O => \N__54453\,
            I => comm_state_3
        );

    \I__13322\ : Odrv4
    port map (
            O => \N__54446\,
            I => comm_state_3
        );

    \I__13321\ : CEMux
    port map (
            O => \N__54431\,
            I => \N__54428\
        );

    \I__13320\ : LocalMux
    port map (
            O => \N__54428\,
            I => \N__54425\
        );

    \I__13319\ : Span4Mux_h
    port map (
            O => \N__54425\,
            I => \N__54422\
        );

    \I__13318\ : Span4Mux_h
    port map (
            O => \N__54422\,
            I => \N__54419\
        );

    \I__13317\ : Odrv4
    port map (
            O => \N__54419\,
            I => n11377
        );

    \I__13316\ : SRMux
    port map (
            O => \N__54416\,
            I => \N__54413\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__54413\,
            I => \N__54410\
        );

    \I__13314\ : Odrv4
    port map (
            O => \N__54410\,
            I => \comm_spi.data_tx_7__N_770\
        );

    \I__13313\ : InMux
    port map (
            O => \N__54407\,
            I => \N__54404\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__54404\,
            I => \N__54401\
        );

    \I__13311\ : Sp12to4
    port map (
            O => \N__54401\,
            I => \N__54398\
        );

    \I__13310\ : Odrv12
    port map (
            O => \N__54398\,
            I => comm_buf_5_6
        );

    \I__13309\ : InMux
    port map (
            O => \N__54395\,
            I => \N__54392\
        );

    \I__13308\ : LocalMux
    port map (
            O => \N__54392\,
            I => \N__54389\
        );

    \I__13307\ : Span12Mux_h
    port map (
            O => \N__54389\,
            I => \N__54386\
        );

    \I__13306\ : Odrv12
    port map (
            O => \N__54386\,
            I => comm_buf_4_6
        );

    \I__13305\ : CascadeMux
    port map (
            O => \N__54383\,
            I => \N__54375\
        );

    \I__13304\ : InMux
    port map (
            O => \N__54382\,
            I => \N__54356\
        );

    \I__13303\ : InMux
    port map (
            O => \N__54381\,
            I => \N__54356\
        );

    \I__13302\ : InMux
    port map (
            O => \N__54380\,
            I => \N__54356\
        );

    \I__13301\ : InMux
    port map (
            O => \N__54379\,
            I => \N__54356\
        );

    \I__13300\ : InMux
    port map (
            O => \N__54378\,
            I => \N__54356\
        );

    \I__13299\ : InMux
    port map (
            O => \N__54375\,
            I => \N__54353\
        );

    \I__13298\ : CascadeMux
    port map (
            O => \N__54374\,
            I => \N__54348\
        );

    \I__13297\ : InMux
    port map (
            O => \N__54373\,
            I => \N__54332\
        );

    \I__13296\ : InMux
    port map (
            O => \N__54372\,
            I => \N__54332\
        );

    \I__13295\ : InMux
    port map (
            O => \N__54371\,
            I => \N__54332\
        );

    \I__13294\ : InMux
    port map (
            O => \N__54370\,
            I => \N__54332\
        );

    \I__13293\ : InMux
    port map (
            O => \N__54369\,
            I => \N__54332\
        );

    \I__13292\ : InMux
    port map (
            O => \N__54368\,
            I => \N__54324\
        );

    \I__13291\ : CascadeMux
    port map (
            O => \N__54367\,
            I => \N__54321\
        );

    \I__13290\ : LocalMux
    port map (
            O => \N__54356\,
            I => \N__54315\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__54353\,
            I => \N__54312\
        );

    \I__13288\ : InMux
    port map (
            O => \N__54352\,
            I => \N__54309\
        );

    \I__13287\ : InMux
    port map (
            O => \N__54351\,
            I => \N__54303\
        );

    \I__13286\ : InMux
    port map (
            O => \N__54348\,
            I => \N__54303\
        );

    \I__13285\ : InMux
    port map (
            O => \N__54347\,
            I => \N__54298\
        );

    \I__13284\ : InMux
    port map (
            O => \N__54346\,
            I => \N__54298\
        );

    \I__13283\ : InMux
    port map (
            O => \N__54345\,
            I => \N__54291\
        );

    \I__13282\ : InMux
    port map (
            O => \N__54344\,
            I => \N__54291\
        );

    \I__13281\ : InMux
    port map (
            O => \N__54343\,
            I => \N__54291\
        );

    \I__13280\ : LocalMux
    port map (
            O => \N__54332\,
            I => \N__54284\
        );

    \I__13279\ : InMux
    port map (
            O => \N__54331\,
            I => \N__54273\
        );

    \I__13278\ : InMux
    port map (
            O => \N__54330\,
            I => \N__54273\
        );

    \I__13277\ : InMux
    port map (
            O => \N__54329\,
            I => \N__54273\
        );

    \I__13276\ : InMux
    port map (
            O => \N__54328\,
            I => \N__54273\
        );

    \I__13275\ : InMux
    port map (
            O => \N__54327\,
            I => \N__54273\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__54324\,
            I => \N__54266\
        );

    \I__13273\ : InMux
    port map (
            O => \N__54321\,
            I => \N__54257\
        );

    \I__13272\ : InMux
    port map (
            O => \N__54320\,
            I => \N__54257\
        );

    \I__13271\ : InMux
    port map (
            O => \N__54319\,
            I => \N__54257\
        );

    \I__13270\ : InMux
    port map (
            O => \N__54318\,
            I => \N__54257\
        );

    \I__13269\ : Span4Mux_v
    port map (
            O => \N__54315\,
            I => \N__54254\
        );

    \I__13268\ : Span4Mux_h
    port map (
            O => \N__54312\,
            I => \N__54249\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54249\
        );

    \I__13266\ : InMux
    port map (
            O => \N__54308\,
            I => \N__54246\
        );

    \I__13265\ : LocalMux
    port map (
            O => \N__54303\,
            I => \N__54239\
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__54298\,
            I => \N__54239\
        );

    \I__13263\ : LocalMux
    port map (
            O => \N__54291\,
            I => \N__54239\
        );

    \I__13262\ : InMux
    port map (
            O => \N__54290\,
            I => \N__54230\
        );

    \I__13261\ : InMux
    port map (
            O => \N__54289\,
            I => \N__54230\
        );

    \I__13260\ : InMux
    port map (
            O => \N__54288\,
            I => \N__54230\
        );

    \I__13259\ : InMux
    port map (
            O => \N__54287\,
            I => \N__54230\
        );

    \I__13258\ : Span4Mux_v
    port map (
            O => \N__54284\,
            I => \N__54225\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__54273\,
            I => \N__54225\
        );

    \I__13256\ : InMux
    port map (
            O => \N__54272\,
            I => \N__54216\
        );

    \I__13255\ : InMux
    port map (
            O => \N__54271\,
            I => \N__54216\
        );

    \I__13254\ : InMux
    port map (
            O => \N__54270\,
            I => \N__54216\
        );

    \I__13253\ : InMux
    port map (
            O => \N__54269\,
            I => \N__54216\
        );

    \I__13252\ : Span4Mux_v
    port map (
            O => \N__54266\,
            I => \N__54207\
        );

    \I__13251\ : LocalMux
    port map (
            O => \N__54257\,
            I => \N__54207\
        );

    \I__13250\ : Span4Mux_h
    port map (
            O => \N__54254\,
            I => \N__54207\
        );

    \I__13249\ : Span4Mux_v
    port map (
            O => \N__54249\,
            I => \N__54207\
        );

    \I__13248\ : LocalMux
    port map (
            O => \N__54246\,
            I => \N__54204\
        );

    \I__13247\ : Odrv4
    port map (
            O => \N__54239\,
            I => comm_index_0
        );

    \I__13246\ : LocalMux
    port map (
            O => \N__54230\,
            I => comm_index_0
        );

    \I__13245\ : Odrv4
    port map (
            O => \N__54225\,
            I => comm_index_0
        );

    \I__13244\ : LocalMux
    port map (
            O => \N__54216\,
            I => comm_index_0
        );

    \I__13243\ : Odrv4
    port map (
            O => \N__54207\,
            I => comm_index_0
        );

    \I__13242\ : Odrv12
    port map (
            O => \N__54204\,
            I => comm_index_0
        );

    \I__13241\ : InMux
    port map (
            O => \N__54191\,
            I => \N__54188\
        );

    \I__13240\ : LocalMux
    port map (
            O => \N__54188\,
            I => \N__54185\
        );

    \I__13239\ : Span4Mux_h
    port map (
            O => \N__54185\,
            I => \N__54182\
        );

    \I__13238\ : Odrv4
    port map (
            O => \N__54182\,
            I => n4_adj_1585
        );

    \I__13237\ : InMux
    port map (
            O => \N__54179\,
            I => \N__54151\
        );

    \I__13236\ : InMux
    port map (
            O => \N__54178\,
            I => \N__54151\
        );

    \I__13235\ : InMux
    port map (
            O => \N__54177\,
            I => \N__54151\
        );

    \I__13234\ : InMux
    port map (
            O => \N__54176\,
            I => \N__54151\
        );

    \I__13233\ : InMux
    port map (
            O => \N__54175\,
            I => \N__54151\
        );

    \I__13232\ : InMux
    port map (
            O => \N__54174\,
            I => \N__54151\
        );

    \I__13231\ : CascadeMux
    port map (
            O => \N__54173\,
            I => \N__54146\
        );

    \I__13230\ : CascadeMux
    port map (
            O => \N__54172\,
            I => \N__54142\
        );

    \I__13229\ : InMux
    port map (
            O => \N__54171\,
            I => \N__54133\
        );

    \I__13228\ : InMux
    port map (
            O => \N__54170\,
            I => \N__54130\
        );

    \I__13227\ : InMux
    port map (
            O => \N__54169\,
            I => \N__54125\
        );

    \I__13226\ : InMux
    port map (
            O => \N__54168\,
            I => \N__54113\
        );

    \I__13225\ : InMux
    port map (
            O => \N__54167\,
            I => \N__54113\
        );

    \I__13224\ : InMux
    port map (
            O => \N__54166\,
            I => \N__54113\
        );

    \I__13223\ : InMux
    port map (
            O => \N__54165\,
            I => \N__54113\
        );

    \I__13222\ : InMux
    port map (
            O => \N__54164\,
            I => \N__54113\
        );

    \I__13221\ : LocalMux
    port map (
            O => \N__54151\,
            I => \N__54110\
        );

    \I__13220\ : InMux
    port map (
            O => \N__54150\,
            I => \N__54107\
        );

    \I__13219\ : InMux
    port map (
            O => \N__54149\,
            I => \N__54095\
        );

    \I__13218\ : InMux
    port map (
            O => \N__54146\,
            I => \N__54095\
        );

    \I__13217\ : InMux
    port map (
            O => \N__54145\,
            I => \N__54095\
        );

    \I__13216\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54095\
        );

    \I__13215\ : InMux
    port map (
            O => \N__54141\,
            I => \N__54095\
        );

    \I__13214\ : CascadeMux
    port map (
            O => \N__54140\,
            I => \N__54092\
        );

    \I__13213\ : InMux
    port map (
            O => \N__54139\,
            I => \N__54064\
        );

    \I__13212\ : InMux
    port map (
            O => \N__54138\,
            I => \N__54057\
        );

    \I__13211\ : InMux
    port map (
            O => \N__54137\,
            I => \N__54057\
        );

    \I__13210\ : InMux
    port map (
            O => \N__54136\,
            I => \N__54057\
        );

    \I__13209\ : LocalMux
    port map (
            O => \N__54133\,
            I => \N__54048\
        );

    \I__13208\ : LocalMux
    port map (
            O => \N__54130\,
            I => \N__54045\
        );

    \I__13207\ : InMux
    port map (
            O => \N__54129\,
            I => \N__54040\
        );

    \I__13206\ : InMux
    port map (
            O => \N__54128\,
            I => \N__54040\
        );

    \I__13205\ : LocalMux
    port map (
            O => \N__54125\,
            I => \N__54037\
        );

    \I__13204\ : InMux
    port map (
            O => \N__54124\,
            I => \N__54023\
        );

    \I__13203\ : LocalMux
    port map (
            O => \N__54113\,
            I => \N__54015\
        );

    \I__13202\ : Span4Mux_h
    port map (
            O => \N__54110\,
            I => \N__54015\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__54107\,
            I => \N__54015\
        );

    \I__13200\ : InMux
    port map (
            O => \N__54106\,
            I => \N__54012\
        );

    \I__13199\ : LocalMux
    port map (
            O => \N__54095\,
            I => \N__54009\
        );

    \I__13198\ : InMux
    port map (
            O => \N__54092\,
            I => \N__53998\
        );

    \I__13197\ : InMux
    port map (
            O => \N__54091\,
            I => \N__53998\
        );

    \I__13196\ : InMux
    port map (
            O => \N__54090\,
            I => \N__53998\
        );

    \I__13195\ : InMux
    port map (
            O => \N__54089\,
            I => \N__53991\
        );

    \I__13194\ : InMux
    port map (
            O => \N__54088\,
            I => \N__53988\
        );

    \I__13193\ : InMux
    port map (
            O => \N__54087\,
            I => \N__53985\
        );

    \I__13192\ : InMux
    port map (
            O => \N__54086\,
            I => \N__53982\
        );

    \I__13191\ : InMux
    port map (
            O => \N__54085\,
            I => \N__53965\
        );

    \I__13190\ : InMux
    port map (
            O => \N__54084\,
            I => \N__53965\
        );

    \I__13189\ : InMux
    port map (
            O => \N__54083\,
            I => \N__53965\
        );

    \I__13188\ : InMux
    port map (
            O => \N__54082\,
            I => \N__53965\
        );

    \I__13187\ : InMux
    port map (
            O => \N__54081\,
            I => \N__53965\
        );

    \I__13186\ : InMux
    port map (
            O => \N__54080\,
            I => \N__53965\
        );

    \I__13185\ : InMux
    port map (
            O => \N__54079\,
            I => \N__53965\
        );

    \I__13184\ : InMux
    port map (
            O => \N__54078\,
            I => \N__53965\
        );

    \I__13183\ : InMux
    port map (
            O => \N__54077\,
            I => \N__53960\
        );

    \I__13182\ : InMux
    port map (
            O => \N__54076\,
            I => \N__53952\
        );

    \I__13181\ : InMux
    port map (
            O => \N__54075\,
            I => \N__53947\
        );

    \I__13180\ : InMux
    port map (
            O => \N__54074\,
            I => \N__53930\
        );

    \I__13179\ : InMux
    port map (
            O => \N__54073\,
            I => \N__53930\
        );

    \I__13178\ : InMux
    port map (
            O => \N__54072\,
            I => \N__53930\
        );

    \I__13177\ : InMux
    port map (
            O => \N__54071\,
            I => \N__53930\
        );

    \I__13176\ : InMux
    port map (
            O => \N__54070\,
            I => \N__53930\
        );

    \I__13175\ : InMux
    port map (
            O => \N__54069\,
            I => \N__53930\
        );

    \I__13174\ : InMux
    port map (
            O => \N__54068\,
            I => \N__53930\
        );

    \I__13173\ : InMux
    port map (
            O => \N__54067\,
            I => \N__53930\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__54064\,
            I => \N__53925\
        );

    \I__13171\ : LocalMux
    port map (
            O => \N__54057\,
            I => \N__53925\
        );

    \I__13170\ : CascadeMux
    port map (
            O => \N__54056\,
            I => \N__53922\
        );

    \I__13169\ : InMux
    port map (
            O => \N__54055\,
            I => \N__53918\
        );

    \I__13168\ : InMux
    port map (
            O => \N__54054\,
            I => \N__53914\
        );

    \I__13167\ : InMux
    port map (
            O => \N__54053\,
            I => \N__53911\
        );

    \I__13166\ : InMux
    port map (
            O => \N__54052\,
            I => \N__53908\
        );

    \I__13165\ : InMux
    port map (
            O => \N__54051\,
            I => \N__53905\
        );

    \I__13164\ : Span4Mux_h
    port map (
            O => \N__54048\,
            I => \N__53902\
        );

    \I__13163\ : Span4Mux_h
    port map (
            O => \N__54045\,
            I => \N__53895\
        );

    \I__13162\ : LocalMux
    port map (
            O => \N__54040\,
            I => \N__53895\
        );

    \I__13161\ : Span4Mux_h
    port map (
            O => \N__54037\,
            I => \N__53895\
        );

    \I__13160\ : InMux
    port map (
            O => \N__54036\,
            I => \N__53892\
        );

    \I__13159\ : InMux
    port map (
            O => \N__54035\,
            I => \N__53885\
        );

    \I__13158\ : InMux
    port map (
            O => \N__54034\,
            I => \N__53885\
        );

    \I__13157\ : InMux
    port map (
            O => \N__54033\,
            I => \N__53885\
        );

    \I__13156\ : InMux
    port map (
            O => \N__54032\,
            I => \N__53878\
        );

    \I__13155\ : InMux
    port map (
            O => \N__54031\,
            I => \N__53878\
        );

    \I__13154\ : InMux
    port map (
            O => \N__54030\,
            I => \N__53878\
        );

    \I__13153\ : InMux
    port map (
            O => \N__54029\,
            I => \N__53875\
        );

    \I__13152\ : InMux
    port map (
            O => \N__54028\,
            I => \N__53872\
        );

    \I__13151\ : InMux
    port map (
            O => \N__54027\,
            I => \N__53869\
        );

    \I__13150\ : InMux
    port map (
            O => \N__54026\,
            I => \N__53866\
        );

    \I__13149\ : LocalMux
    port map (
            O => \N__54023\,
            I => \N__53863\
        );

    \I__13148\ : InMux
    port map (
            O => \N__54022\,
            I => \N__53859\
        );

    \I__13147\ : Span4Mux_v
    port map (
            O => \N__54015\,
            I => \N__53856\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__54012\,
            I => \N__53851\
        );

    \I__13145\ : Span4Mux_v
    port map (
            O => \N__54009\,
            I => \N__53851\
        );

    \I__13144\ : InMux
    port map (
            O => \N__54008\,
            I => \N__53844\
        );

    \I__13143\ : InMux
    port map (
            O => \N__54007\,
            I => \N__53844\
        );

    \I__13142\ : InMux
    port map (
            O => \N__54006\,
            I => \N__53844\
        );

    \I__13141\ : InMux
    port map (
            O => \N__54005\,
            I => \N__53839\
        );

    \I__13140\ : LocalMux
    port map (
            O => \N__53998\,
            I => \N__53836\
        );

    \I__13139\ : InMux
    port map (
            O => \N__53997\,
            I => \N__53829\
        );

    \I__13138\ : InMux
    port map (
            O => \N__53996\,
            I => \N__53829\
        );

    \I__13137\ : InMux
    port map (
            O => \N__53995\,
            I => \N__53829\
        );

    \I__13136\ : InMux
    port map (
            O => \N__53994\,
            I => \N__53826\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__53991\,
            I => \N__53817\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__53988\,
            I => \N__53817\
        );

    \I__13133\ : LocalMux
    port map (
            O => \N__53985\,
            I => \N__53817\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__53982\,
            I => \N__53817\
        );

    \I__13131\ : LocalMux
    port map (
            O => \N__53965\,
            I => \N__53814\
        );

    \I__13130\ : InMux
    port map (
            O => \N__53964\,
            I => \N__53807\
        );

    \I__13129\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53807\
        );

    \I__13128\ : LocalMux
    port map (
            O => \N__53960\,
            I => \N__53801\
        );

    \I__13127\ : InMux
    port map (
            O => \N__53959\,
            I => \N__53794\
        );

    \I__13126\ : InMux
    port map (
            O => \N__53958\,
            I => \N__53794\
        );

    \I__13125\ : InMux
    port map (
            O => \N__53957\,
            I => \N__53794\
        );

    \I__13124\ : InMux
    port map (
            O => \N__53956\,
            I => \N__53789\
        );

    \I__13123\ : InMux
    port map (
            O => \N__53955\,
            I => \N__53789\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__53952\,
            I => \N__53783\
        );

    \I__13121\ : InMux
    port map (
            O => \N__53951\,
            I => \N__53778\
        );

    \I__13120\ : InMux
    port map (
            O => \N__53950\,
            I => \N__53778\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__53947\,
            I => \N__53775\
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__53930\,
            I => \N__53765\
        );

    \I__13117\ : Span4Mux_v
    port map (
            O => \N__53925\,
            I => \N__53765\
        );

    \I__13116\ : InMux
    port map (
            O => \N__53922\,
            I => \N__53760\
        );

    \I__13115\ : InMux
    port map (
            O => \N__53921\,
            I => \N__53760\
        );

    \I__13114\ : LocalMux
    port map (
            O => \N__53918\,
            I => \N__53757\
        );

    \I__13113\ : InMux
    port map (
            O => \N__53917\,
            I => \N__53754\
        );

    \I__13112\ : LocalMux
    port map (
            O => \N__53914\,
            I => \N__53741\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__53911\,
            I => \N__53741\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__53908\,
            I => \N__53741\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53741\
        );

    \I__13108\ : Span4Mux_h
    port map (
            O => \N__53902\,
            I => \N__53741\
        );

    \I__13107\ : Span4Mux_v
    port map (
            O => \N__53895\,
            I => \N__53741\
        );

    \I__13106\ : LocalMux
    port map (
            O => \N__53892\,
            I => \N__53732\
        );

    \I__13105\ : LocalMux
    port map (
            O => \N__53885\,
            I => \N__53732\
        );

    \I__13104\ : LocalMux
    port map (
            O => \N__53878\,
            I => \N__53732\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__53875\,
            I => \N__53732\
        );

    \I__13102\ : LocalMux
    port map (
            O => \N__53872\,
            I => \N__53729\
        );

    \I__13101\ : LocalMux
    port map (
            O => \N__53869\,
            I => \N__53722\
        );

    \I__13100\ : LocalMux
    port map (
            O => \N__53866\,
            I => \N__53722\
        );

    \I__13099\ : Span4Mux_h
    port map (
            O => \N__53863\,
            I => \N__53722\
        );

    \I__13098\ : InMux
    port map (
            O => \N__53862\,
            I => \N__53719\
        );

    \I__13097\ : LocalMux
    port map (
            O => \N__53859\,
            I => \N__53710\
        );

    \I__13096\ : Span4Mux_h
    port map (
            O => \N__53856\,
            I => \N__53710\
        );

    \I__13095\ : Span4Mux_h
    port map (
            O => \N__53851\,
            I => \N__53710\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__53844\,
            I => \N__53710\
        );

    \I__13093\ : InMux
    port map (
            O => \N__53843\,
            I => \N__53705\
        );

    \I__13092\ : InMux
    port map (
            O => \N__53842\,
            I => \N__53705\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__53839\,
            I => \N__53698\
        );

    \I__13090\ : Sp12to4
    port map (
            O => \N__53836\,
            I => \N__53698\
        );

    \I__13089\ : LocalMux
    port map (
            O => \N__53829\,
            I => \N__53698\
        );

    \I__13088\ : LocalMux
    port map (
            O => \N__53826\,
            I => \N__53691\
        );

    \I__13087\ : Span4Mux_v
    port map (
            O => \N__53817\,
            I => \N__53691\
        );

    \I__13086\ : Span4Mux_v
    port map (
            O => \N__53814\,
            I => \N__53691\
        );

    \I__13085\ : InMux
    port map (
            O => \N__53813\,
            I => \N__53686\
        );

    \I__13084\ : InMux
    port map (
            O => \N__53812\,
            I => \N__53686\
        );

    \I__13083\ : LocalMux
    port map (
            O => \N__53807\,
            I => \N__53683\
        );

    \I__13082\ : InMux
    port map (
            O => \N__53806\,
            I => \N__53676\
        );

    \I__13081\ : InMux
    port map (
            O => \N__53805\,
            I => \N__53676\
        );

    \I__13080\ : InMux
    port map (
            O => \N__53804\,
            I => \N__53676\
        );

    \I__13079\ : Span4Mux_h
    port map (
            O => \N__53801\,
            I => \N__53669\
        );

    \I__13078\ : LocalMux
    port map (
            O => \N__53794\,
            I => \N__53669\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__53789\,
            I => \N__53669\
        );

    \I__13076\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53662\
        );

    \I__13075\ : InMux
    port map (
            O => \N__53787\,
            I => \N__53662\
        );

    \I__13074\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53662\
        );

    \I__13073\ : Span4Mux_v
    port map (
            O => \N__53783\,
            I => \N__53655\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__53778\,
            I => \N__53655\
        );

    \I__13071\ : Span4Mux_h
    port map (
            O => \N__53775\,
            I => \N__53655\
        );

    \I__13070\ : InMux
    port map (
            O => \N__53774\,
            I => \N__53650\
        );

    \I__13069\ : InMux
    port map (
            O => \N__53773\,
            I => \N__53650\
        );

    \I__13068\ : InMux
    port map (
            O => \N__53772\,
            I => \N__53643\
        );

    \I__13067\ : InMux
    port map (
            O => \N__53771\,
            I => \N__53643\
        );

    \I__13066\ : InMux
    port map (
            O => \N__53770\,
            I => \N__53643\
        );

    \I__13065\ : Span4Mux_h
    port map (
            O => \N__53765\,
            I => \N__53628\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__53760\,
            I => \N__53628\
        );

    \I__13063\ : Span4Mux_v
    port map (
            O => \N__53757\,
            I => \N__53628\
        );

    \I__13062\ : LocalMux
    port map (
            O => \N__53754\,
            I => \N__53628\
        );

    \I__13061\ : Span4Mux_v
    port map (
            O => \N__53741\,
            I => \N__53628\
        );

    \I__13060\ : Span4Mux_v
    port map (
            O => \N__53732\,
            I => \N__53628\
        );

    \I__13059\ : Span4Mux_v
    port map (
            O => \N__53729\,
            I => \N__53628\
        );

    \I__13058\ : Span4Mux_v
    port map (
            O => \N__53722\,
            I => \N__53621\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__53719\,
            I => \N__53621\
        );

    \I__13056\ : Span4Mux_h
    port map (
            O => \N__53710\,
            I => \N__53621\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__53705\,
            I => \N__53616\
        );

    \I__13054\ : Span12Mux_v
    port map (
            O => \N__53698\,
            I => \N__53616\
        );

    \I__13053\ : Odrv4
    port map (
            O => \N__53691\,
            I => comm_state_1
        );

    \I__13052\ : LocalMux
    port map (
            O => \N__53686\,
            I => comm_state_1
        );

    \I__13051\ : Odrv4
    port map (
            O => \N__53683\,
            I => comm_state_1
        );

    \I__13050\ : LocalMux
    port map (
            O => \N__53676\,
            I => comm_state_1
        );

    \I__13049\ : Odrv4
    port map (
            O => \N__53669\,
            I => comm_state_1
        );

    \I__13048\ : LocalMux
    port map (
            O => \N__53662\,
            I => comm_state_1
        );

    \I__13047\ : Odrv4
    port map (
            O => \N__53655\,
            I => comm_state_1
        );

    \I__13046\ : LocalMux
    port map (
            O => \N__53650\,
            I => comm_state_1
        );

    \I__13045\ : LocalMux
    port map (
            O => \N__53643\,
            I => comm_state_1
        );

    \I__13044\ : Odrv4
    port map (
            O => \N__53628\,
            I => comm_state_1
        );

    \I__13043\ : Odrv4
    port map (
            O => \N__53621\,
            I => comm_state_1
        );

    \I__13042\ : Odrv12
    port map (
            O => \N__53616\,
            I => comm_state_1
        );

    \I__13041\ : InMux
    port map (
            O => \N__53591\,
            I => \N__53583\
        );

    \I__13040\ : InMux
    port map (
            O => \N__53590\,
            I => \N__53572\
        );

    \I__13039\ : InMux
    port map (
            O => \N__53589\,
            I => \N__53572\
        );

    \I__13038\ : InMux
    port map (
            O => \N__53588\,
            I => \N__53572\
        );

    \I__13037\ : InMux
    port map (
            O => \N__53587\,
            I => \N__53572\
        );

    \I__13036\ : InMux
    port map (
            O => \N__53586\,
            I => \N__53569\
        );

    \I__13035\ : LocalMux
    port map (
            O => \N__53583\,
            I => \N__53558\
        );

    \I__13034\ : InMux
    port map (
            O => \N__53582\,
            I => \N__53555\
        );

    \I__13033\ : InMux
    port map (
            O => \N__53581\,
            I => \N__53550\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__53572\,
            I => \N__53545\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__53569\,
            I => \N__53542\
        );

    \I__13030\ : InMux
    port map (
            O => \N__53568\,
            I => \N__53539\
        );

    \I__13029\ : InMux
    port map (
            O => \N__53567\,
            I => \N__53534\
        );

    \I__13028\ : InMux
    port map (
            O => \N__53566\,
            I => \N__53531\
        );

    \I__13027\ : InMux
    port map (
            O => \N__53565\,
            I => \N__53524\
        );

    \I__13026\ : InMux
    port map (
            O => \N__53564\,
            I => \N__53524\
        );

    \I__13025\ : InMux
    port map (
            O => \N__53563\,
            I => \N__53524\
        );

    \I__13024\ : InMux
    port map (
            O => \N__53562\,
            I => \N__53521\
        );

    \I__13023\ : InMux
    port map (
            O => \N__53561\,
            I => \N__53513\
        );

    \I__13022\ : Span4Mux_v
    port map (
            O => \N__53558\,
            I => \N__53510\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__53555\,
            I => \N__53507\
        );

    \I__13020\ : InMux
    port map (
            O => \N__53554\,
            I => \N__53498\
        );

    \I__13019\ : InMux
    port map (
            O => \N__53553\,
            I => \N__53498\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__53550\,
            I => \N__53492\
        );

    \I__13017\ : InMux
    port map (
            O => \N__53549\,
            I => \N__53489\
        );

    \I__13016\ : InMux
    port map (
            O => \N__53548\,
            I => \N__53486\
        );

    \I__13015\ : Span4Mux_v
    port map (
            O => \N__53545\,
            I => \N__53479\
        );

    \I__13014\ : Span4Mux_v
    port map (
            O => \N__53542\,
            I => \N__53479\
        );

    \I__13013\ : LocalMux
    port map (
            O => \N__53539\,
            I => \N__53479\
        );

    \I__13012\ : InMux
    port map (
            O => \N__53538\,
            I => \N__53474\
        );

    \I__13011\ : InMux
    port map (
            O => \N__53537\,
            I => \N__53474\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__53534\,
            I => \N__53471\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__53531\,
            I => \N__53468\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__53524\,
            I => \N__53460\
        );

    \I__13007\ : LocalMux
    port map (
            O => \N__53521\,
            I => \N__53460\
        );

    \I__13006\ : InMux
    port map (
            O => \N__53520\,
            I => \N__53455\
        );

    \I__13005\ : InMux
    port map (
            O => \N__53519\,
            I => \N__53455\
        );

    \I__13004\ : InMux
    port map (
            O => \N__53518\,
            I => \N__53448\
        );

    \I__13003\ : InMux
    port map (
            O => \N__53517\,
            I => \N__53448\
        );

    \I__13002\ : InMux
    port map (
            O => \N__53516\,
            I => \N__53448\
        );

    \I__13001\ : LocalMux
    port map (
            O => \N__53513\,
            I => \N__53443\
        );

    \I__13000\ : Span4Mux_h
    port map (
            O => \N__53510\,
            I => \N__53443\
        );

    \I__12999\ : Span4Mux_v
    port map (
            O => \N__53507\,
            I => \N__53440\
        );

    \I__12998\ : InMux
    port map (
            O => \N__53506\,
            I => \N__53435\
        );

    \I__12997\ : InMux
    port map (
            O => \N__53505\,
            I => \N__53435\
        );

    \I__12996\ : InMux
    port map (
            O => \N__53504\,
            I => \N__53430\
        );

    \I__12995\ : InMux
    port map (
            O => \N__53503\,
            I => \N__53430\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__53498\,
            I => \N__53427\
        );

    \I__12993\ : InMux
    port map (
            O => \N__53497\,
            I => \N__53420\
        );

    \I__12992\ : InMux
    port map (
            O => \N__53496\,
            I => \N__53420\
        );

    \I__12991\ : InMux
    port map (
            O => \N__53495\,
            I => \N__53420\
        );

    \I__12990\ : Span4Mux_v
    port map (
            O => \N__53492\,
            I => \N__53417\
        );

    \I__12989\ : LocalMux
    port map (
            O => \N__53489\,
            I => \N__53414\
        );

    \I__12988\ : LocalMux
    port map (
            O => \N__53486\,
            I => \N__53411\
        );

    \I__12987\ : Span4Mux_v
    port map (
            O => \N__53479\,
            I => \N__53408\
        );

    \I__12986\ : LocalMux
    port map (
            O => \N__53474\,
            I => \N__53405\
        );

    \I__12985\ : Span4Mux_v
    port map (
            O => \N__53471\,
            I => \N__53400\
        );

    \I__12984\ : Span4Mux_v
    port map (
            O => \N__53468\,
            I => \N__53400\
        );

    \I__12983\ : InMux
    port map (
            O => \N__53467\,
            I => \N__53393\
        );

    \I__12982\ : InMux
    port map (
            O => \N__53466\,
            I => \N__53393\
        );

    \I__12981\ : InMux
    port map (
            O => \N__53465\,
            I => \N__53393\
        );

    \I__12980\ : Span4Mux_h
    port map (
            O => \N__53460\,
            I => \N__53386\
        );

    \I__12979\ : LocalMux
    port map (
            O => \N__53455\,
            I => \N__53386\
        );

    \I__12978\ : LocalMux
    port map (
            O => \N__53448\,
            I => \N__53386\
        );

    \I__12977\ : Span4Mux_h
    port map (
            O => \N__53443\,
            I => \N__53383\
        );

    \I__12976\ : Span4Mux_v
    port map (
            O => \N__53440\,
            I => \N__53364\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__53435\,
            I => \N__53364\
        );

    \I__12974\ : LocalMux
    port map (
            O => \N__53430\,
            I => \N__53364\
        );

    \I__12973\ : Span4Mux_v
    port map (
            O => \N__53427\,
            I => \N__53364\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__53420\,
            I => \N__53364\
        );

    \I__12971\ : Span4Mux_v
    port map (
            O => \N__53417\,
            I => \N__53364\
        );

    \I__12970\ : Span4Mux_v
    port map (
            O => \N__53414\,
            I => \N__53364\
        );

    \I__12969\ : Span4Mux_v
    port map (
            O => \N__53411\,
            I => \N__53364\
        );

    \I__12968\ : Span4Mux_h
    port map (
            O => \N__53408\,
            I => \N__53364\
        );

    \I__12967\ : Odrv4
    port map (
            O => \N__53405\,
            I => comm_state_0
        );

    \I__12966\ : Odrv4
    port map (
            O => \N__53400\,
            I => comm_state_0
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__53393\,
            I => comm_state_0
        );

    \I__12964\ : Odrv4
    port map (
            O => \N__53386\,
            I => comm_state_0
        );

    \I__12963\ : Odrv4
    port map (
            O => \N__53383\,
            I => comm_state_0
        );

    \I__12962\ : Odrv4
    port map (
            O => \N__53364\,
            I => comm_state_0
        );

    \I__12961\ : CascadeMux
    port map (
            O => \N__53351\,
            I => \N__53347\
        );

    \I__12960\ : InMux
    port map (
            O => \N__53350\,
            I => \N__53341\
        );

    \I__12959\ : InMux
    port map (
            O => \N__53347\,
            I => \N__53341\
        );

    \I__12958\ : InMux
    port map (
            O => \N__53346\,
            I => \N__53338\
        );

    \I__12957\ : LocalMux
    port map (
            O => \N__53341\,
            I => \N__53333\
        );

    \I__12956\ : LocalMux
    port map (
            O => \N__53338\,
            I => \N__53333\
        );

    \I__12955\ : Span4Mux_h
    port map (
            O => \N__53333\,
            I => \N__53330\
        );

    \I__12954\ : Odrv4
    port map (
            O => \N__53330\,
            I => n9270
        );

    \I__12953\ : InMux
    port map (
            O => \N__53327\,
            I => \N__53321\
        );

    \I__12952\ : InMux
    port map (
            O => \N__53326\,
            I => \N__53318\
        );

    \I__12951\ : InMux
    port map (
            O => \N__53325\,
            I => \N__53313\
        );

    \I__12950\ : InMux
    port map (
            O => \N__53324\,
            I => \N__53313\
        );

    \I__12949\ : LocalMux
    port map (
            O => \N__53321\,
            I => \comm_spi.n22670\
        );

    \I__12948\ : LocalMux
    port map (
            O => \N__53318\,
            I => \comm_spi.n22670\
        );

    \I__12947\ : LocalMux
    port map (
            O => \N__53313\,
            I => \comm_spi.n22670\
        );

    \I__12946\ : InMux
    port map (
            O => \N__53306\,
            I => \N__53303\
        );

    \I__12945\ : LocalMux
    port map (
            O => \N__53303\,
            I => \comm_spi.n14631\
        );

    \I__12944\ : InMux
    port map (
            O => \N__53300\,
            I => \N__53297\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__53297\,
            I => \N__53292\
        );

    \I__12942\ : InMux
    port map (
            O => \N__53296\,
            I => \N__53289\
        );

    \I__12941\ : InMux
    port map (
            O => \N__53295\,
            I => \N__53286\
        );

    \I__12940\ : Odrv4
    port map (
            O => \N__53292\,
            I => \comm_spi.n14616\
        );

    \I__12939\ : LocalMux
    port map (
            O => \N__53289\,
            I => \comm_spi.n14616\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__53286\,
            I => \comm_spi.n14616\
        );

    \I__12937\ : InMux
    port map (
            O => \N__53279\,
            I => \N__53274\
        );

    \I__12936\ : InMux
    port map (
            O => \N__53278\,
            I => \N__53271\
        );

    \I__12935\ : InMux
    port map (
            O => \N__53277\,
            I => \N__53268\
        );

    \I__12934\ : LocalMux
    port map (
            O => \N__53274\,
            I => \N__53265\
        );

    \I__12933\ : LocalMux
    port map (
            O => \N__53271\,
            I => \N__53260\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__53268\,
            I => \N__53260\
        );

    \I__12931\ : Odrv4
    port map (
            O => \N__53265\,
            I => \comm_spi.n14617\
        );

    \I__12930\ : Odrv4
    port map (
            O => \N__53260\,
            I => \comm_spi.n14617\
        );

    \I__12929\ : CascadeMux
    port map (
            O => \N__53255\,
            I => \N__53251\
        );

    \I__12928\ : InMux
    port map (
            O => \N__53254\,
            I => \N__53247\
        );

    \I__12927\ : InMux
    port map (
            O => \N__53251\,
            I => \N__53242\
        );

    \I__12926\ : InMux
    port map (
            O => \N__53250\,
            I => \N__53242\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__53247\,
            I => cmd_rdadctmp_19_adj_1431
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__53242\,
            I => cmd_rdadctmp_19_adj_1431
        );

    \I__12923\ : InMux
    port map (
            O => \N__53237\,
            I => \N__53234\
        );

    \I__12922\ : LocalMux
    port map (
            O => \N__53234\,
            I => \N__53231\
        );

    \I__12921\ : Span4Mux_v
    port map (
            O => \N__53231\,
            I => \N__53226\
        );

    \I__12920\ : InMux
    port map (
            O => \N__53230\,
            I => \N__53223\
        );

    \I__12919\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53220\
        );

    \I__12918\ : Span4Mux_h
    port map (
            O => \N__53226\,
            I => \N__53217\
        );

    \I__12917\ : LocalMux
    port map (
            O => \N__53223\,
            I => \N__53214\
        );

    \I__12916\ : LocalMux
    port map (
            O => \N__53220\,
            I => buf_adcdata_iac_11
        );

    \I__12915\ : Odrv4
    port map (
            O => \N__53217\,
            I => buf_adcdata_iac_11
        );

    \I__12914\ : Odrv12
    port map (
            O => \N__53214\,
            I => buf_adcdata_iac_11
        );

    \I__12913\ : InMux
    port map (
            O => \N__53207\,
            I => \N__53201\
        );

    \I__12912\ : InMux
    port map (
            O => \N__53206\,
            I => \N__53201\
        );

    \I__12911\ : LocalMux
    port map (
            O => \N__53201\,
            I => \N__53195\
        );

    \I__12910\ : InMux
    port map (
            O => \N__53200\,
            I => \N__53192\
        );

    \I__12909\ : InMux
    port map (
            O => \N__53199\,
            I => \N__53189\
        );

    \I__12908\ : InMux
    port map (
            O => \N__53198\,
            I => \N__53186\
        );

    \I__12907\ : Span4Mux_h
    port map (
            O => \N__53195\,
            I => \N__53180\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__53192\,
            I => \N__53172\
        );

    \I__12905\ : LocalMux
    port map (
            O => \N__53189\,
            I => \N__53167\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__53186\,
            I => \N__53167\
        );

    \I__12903\ : InMux
    port map (
            O => \N__53185\,
            I => \N__53163\
        );

    \I__12902\ : InMux
    port map (
            O => \N__53184\,
            I => \N__53160\
        );

    \I__12901\ : InMux
    port map (
            O => \N__53183\,
            I => \N__53157\
        );

    \I__12900\ : Span4Mux_h
    port map (
            O => \N__53180\,
            I => \N__53153\
        );

    \I__12899\ : InMux
    port map (
            O => \N__53179\,
            I => \N__53146\
        );

    \I__12898\ : InMux
    port map (
            O => \N__53178\,
            I => \N__53146\
        );

    \I__12897\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53146\
        );

    \I__12896\ : InMux
    port map (
            O => \N__53176\,
            I => \N__53143\
        );

    \I__12895\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53140\
        );

    \I__12894\ : Span4Mux_h
    port map (
            O => \N__53172\,
            I => \N__53135\
        );

    \I__12893\ : Span4Mux_v
    port map (
            O => \N__53167\,
            I => \N__53135\
        );

    \I__12892\ : InMux
    port map (
            O => \N__53166\,
            I => \N__53132\
        );

    \I__12891\ : LocalMux
    port map (
            O => \N__53163\,
            I => \N__53124\
        );

    \I__12890\ : LocalMux
    port map (
            O => \N__53160\,
            I => \N__53121\
        );

    \I__12889\ : LocalMux
    port map (
            O => \N__53157\,
            I => \N__53118\
        );

    \I__12888\ : CascadeMux
    port map (
            O => \N__53156\,
            I => \N__53113\
        );

    \I__12887\ : Sp12to4
    port map (
            O => \N__53153\,
            I => \N__53110\
        );

    \I__12886\ : LocalMux
    port map (
            O => \N__53146\,
            I => \N__53105\
        );

    \I__12885\ : LocalMux
    port map (
            O => \N__53143\,
            I => \N__53105\
        );

    \I__12884\ : LocalMux
    port map (
            O => \N__53140\,
            I => \N__53102\
        );

    \I__12883\ : Span4Mux_v
    port map (
            O => \N__53135\,
            I => \N__53097\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__53132\,
            I => \N__53097\
        );

    \I__12881\ : InMux
    port map (
            O => \N__53131\,
            I => \N__53092\
        );

    \I__12880\ : InMux
    port map (
            O => \N__53130\,
            I => \N__53092\
        );

    \I__12879\ : InMux
    port map (
            O => \N__53129\,
            I => \N__53085\
        );

    \I__12878\ : InMux
    port map (
            O => \N__53128\,
            I => \N__53085\
        );

    \I__12877\ : InMux
    port map (
            O => \N__53127\,
            I => \N__53085\
        );

    \I__12876\ : Span4Mux_v
    port map (
            O => \N__53124\,
            I => \N__53080\
        );

    \I__12875\ : Span4Mux_v
    port map (
            O => \N__53121\,
            I => \N__53080\
        );

    \I__12874\ : Span4Mux_v
    port map (
            O => \N__53118\,
            I => \N__53077\
        );

    \I__12873\ : InMux
    port map (
            O => \N__53117\,
            I => \N__53070\
        );

    \I__12872\ : InMux
    port map (
            O => \N__53116\,
            I => \N__53070\
        );

    \I__12871\ : InMux
    port map (
            O => \N__53113\,
            I => \N__53070\
        );

    \I__12870\ : Span12Mux_v
    port map (
            O => \N__53110\,
            I => \N__53063\
        );

    \I__12869\ : Span12Mux_v
    port map (
            O => \N__53105\,
            I => \N__53063\
        );

    \I__12868\ : Span4Mux_h
    port map (
            O => \N__53102\,
            I => \N__53060\
        );

    \I__12867\ : Span4Mux_v
    port map (
            O => \N__53097\,
            I => \N__53053\
        );

    \I__12866\ : LocalMux
    port map (
            O => \N__53092\,
            I => \N__53053\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__53085\,
            I => \N__53053\
        );

    \I__12864\ : Span4Mux_v
    port map (
            O => \N__53080\,
            I => \N__53050\
        );

    \I__12863\ : Span4Mux_v
    port map (
            O => \N__53077\,
            I => \N__53047\
        );

    \I__12862\ : LocalMux
    port map (
            O => \N__53070\,
            I => \N__53044\
        );

    \I__12861\ : InMux
    port map (
            O => \N__53069\,
            I => \N__53039\
        );

    \I__12860\ : InMux
    port map (
            O => \N__53068\,
            I => \N__53039\
        );

    \I__12859\ : Span12Mux_h
    port map (
            O => \N__53063\,
            I => \N__53036\
        );

    \I__12858\ : Span4Mux_h
    port map (
            O => \N__53060\,
            I => \N__53033\
        );

    \I__12857\ : Span4Mux_h
    port map (
            O => \N__53053\,
            I => \N__53030\
        );

    \I__12856\ : Span4Mux_v
    port map (
            O => \N__53050\,
            I => \N__53021\
        );

    \I__12855\ : Span4Mux_h
    port map (
            O => \N__53047\,
            I => \N__53021\
        );

    \I__12854\ : Span4Mux_h
    port map (
            O => \N__53044\,
            I => \N__53021\
        );

    \I__12853\ : LocalMux
    port map (
            O => \N__53039\,
            I => \N__53021\
        );

    \I__12852\ : Odrv12
    port map (
            O => \N__53036\,
            I => n20584
        );

    \I__12851\ : Odrv4
    port map (
            O => \N__53033\,
            I => n20584
        );

    \I__12850\ : Odrv4
    port map (
            O => \N__53030\,
            I => n20584
        );

    \I__12849\ : Odrv4
    port map (
            O => \N__53021\,
            I => n20584
        );

    \I__12848\ : InMux
    port map (
            O => \N__53012\,
            I => \N__53008\
        );

    \I__12847\ : InMux
    port map (
            O => \N__53011\,
            I => \N__52986\
        );

    \I__12846\ : LocalMux
    port map (
            O => \N__53008\,
            I => \N__52983\
        );

    \I__12845\ : InMux
    port map (
            O => \N__53007\,
            I => \N__52970\
        );

    \I__12844\ : InMux
    port map (
            O => \N__53006\,
            I => \N__52970\
        );

    \I__12843\ : InMux
    port map (
            O => \N__53005\,
            I => \N__52970\
        );

    \I__12842\ : InMux
    port map (
            O => \N__53004\,
            I => \N__52970\
        );

    \I__12841\ : InMux
    port map (
            O => \N__53003\,
            I => \N__52970\
        );

    \I__12840\ : InMux
    port map (
            O => \N__53002\,
            I => \N__52970\
        );

    \I__12839\ : CascadeMux
    port map (
            O => \N__53001\,
            I => \N__52967\
        );

    \I__12838\ : InMux
    port map (
            O => \N__53000\,
            I => \N__52960\
        );

    \I__12837\ : InMux
    port map (
            O => \N__52999\,
            I => \N__52960\
        );

    \I__12836\ : InMux
    port map (
            O => \N__52998\,
            I => \N__52960\
        );

    \I__12835\ : CascadeMux
    port map (
            O => \N__52997\,
            I => \N__52955\
        );

    \I__12834\ : InMux
    port map (
            O => \N__52996\,
            I => \N__52948\
        );

    \I__12833\ : InMux
    port map (
            O => \N__52995\,
            I => \N__52945\
        );

    \I__12832\ : InMux
    port map (
            O => \N__52994\,
            I => \N__52942\
        );

    \I__12831\ : InMux
    port map (
            O => \N__52993\,
            I => \N__52937\
        );

    \I__12830\ : InMux
    port map (
            O => \N__52992\,
            I => \N__52937\
        );

    \I__12829\ : InMux
    port map (
            O => \N__52991\,
            I => \N__52930\
        );

    \I__12828\ : InMux
    port map (
            O => \N__52990\,
            I => \N__52927\
        );

    \I__12827\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52924\
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__52986\,
            I => \N__52917\
        );

    \I__12825\ : Span4Mux_h
    port map (
            O => \N__52983\,
            I => \N__52917\
        );

    \I__12824\ : LocalMux
    port map (
            O => \N__52970\,
            I => \N__52917\
        );

    \I__12823\ : InMux
    port map (
            O => \N__52967\,
            I => \N__52912\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__52960\,
            I => \N__52908\
        );

    \I__12821\ : InMux
    port map (
            O => \N__52959\,
            I => \N__52903\
        );

    \I__12820\ : InMux
    port map (
            O => \N__52958\,
            I => \N__52903\
        );

    \I__12819\ : InMux
    port map (
            O => \N__52955\,
            I => \N__52900\
        );

    \I__12818\ : InMux
    port map (
            O => \N__52954\,
            I => \N__52891\
        );

    \I__12817\ : InMux
    port map (
            O => \N__52953\,
            I => \N__52891\
        );

    \I__12816\ : InMux
    port map (
            O => \N__52952\,
            I => \N__52891\
        );

    \I__12815\ : InMux
    port map (
            O => \N__52951\,
            I => \N__52891\
        );

    \I__12814\ : LocalMux
    port map (
            O => \N__52948\,
            I => \N__52886\
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__52945\,
            I => \N__52886\
        );

    \I__12812\ : LocalMux
    port map (
            O => \N__52942\,
            I => \N__52881\
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__52937\,
            I => \N__52881\
        );

    \I__12810\ : InMux
    port map (
            O => \N__52936\,
            I => \N__52866\
        );

    \I__12809\ : InMux
    port map (
            O => \N__52935\,
            I => \N__52866\
        );

    \I__12808\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52866\
        );

    \I__12807\ : InMux
    port map (
            O => \N__52933\,
            I => \N__52866\
        );

    \I__12806\ : LocalMux
    port map (
            O => \N__52930\,
            I => \N__52863\
        );

    \I__12805\ : LocalMux
    port map (
            O => \N__52927\,
            I => \N__52858\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__52924\,
            I => \N__52858\
        );

    \I__12803\ : Span4Mux_v
    port map (
            O => \N__52917\,
            I => \N__52855\
        );

    \I__12802\ : CascadeMux
    port map (
            O => \N__52916\,
            I => \N__52851\
        );

    \I__12801\ : InMux
    port map (
            O => \N__52915\,
            I => \N__52841\
        );

    \I__12800\ : LocalMux
    port map (
            O => \N__52912\,
            I => \N__52838\
        );

    \I__12799\ : InMux
    port map (
            O => \N__52911\,
            I => \N__52835\
        );

    \I__12798\ : Span4Mux_h
    port map (
            O => \N__52908\,
            I => \N__52832\
        );

    \I__12797\ : LocalMux
    port map (
            O => \N__52903\,
            I => \N__52829\
        );

    \I__12796\ : LocalMux
    port map (
            O => \N__52900\,
            I => \N__52820\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__52891\,
            I => \N__52820\
        );

    \I__12794\ : Span4Mux_h
    port map (
            O => \N__52886\,
            I => \N__52820\
        );

    \I__12793\ : Span4Mux_h
    port map (
            O => \N__52881\,
            I => \N__52820\
        );

    \I__12792\ : InMux
    port map (
            O => \N__52880\,
            I => \N__52806\
        );

    \I__12791\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52806\
        );

    \I__12790\ : InMux
    port map (
            O => \N__52878\,
            I => \N__52806\
        );

    \I__12789\ : InMux
    port map (
            O => \N__52877\,
            I => \N__52806\
        );

    \I__12788\ : InMux
    port map (
            O => \N__52876\,
            I => \N__52806\
        );

    \I__12787\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52806\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__52866\,
            I => \N__52801\
        );

    \I__12785\ : Span4Mux_v
    port map (
            O => \N__52863\,
            I => \N__52801\
        );

    \I__12784\ : Span4Mux_v
    port map (
            O => \N__52858\,
            I => \N__52796\
        );

    \I__12783\ : Span4Mux_h
    port map (
            O => \N__52855\,
            I => \N__52796\
        );

    \I__12782\ : InMux
    port map (
            O => \N__52854\,
            I => \N__52793\
        );

    \I__12781\ : InMux
    port map (
            O => \N__52851\,
            I => \N__52788\
        );

    \I__12780\ : InMux
    port map (
            O => \N__52850\,
            I => \N__52788\
        );

    \I__12779\ : InMux
    port map (
            O => \N__52849\,
            I => \N__52779\
        );

    \I__12778\ : InMux
    port map (
            O => \N__52848\,
            I => \N__52779\
        );

    \I__12777\ : InMux
    port map (
            O => \N__52847\,
            I => \N__52779\
        );

    \I__12776\ : InMux
    port map (
            O => \N__52846\,
            I => \N__52779\
        );

    \I__12775\ : InMux
    port map (
            O => \N__52845\,
            I => \N__52774\
        );

    \I__12774\ : InMux
    port map (
            O => \N__52844\,
            I => \N__52774\
        );

    \I__12773\ : LocalMux
    port map (
            O => \N__52841\,
            I => \N__52769\
        );

    \I__12772\ : Span4Mux_v
    port map (
            O => \N__52838\,
            I => \N__52769\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__52835\,
            I => \N__52764\
        );

    \I__12770\ : Span4Mux_v
    port map (
            O => \N__52832\,
            I => \N__52764\
        );

    \I__12769\ : Span4Mux_h
    port map (
            O => \N__52829\,
            I => \N__52759\
        );

    \I__12768\ : Span4Mux_v
    port map (
            O => \N__52820\,
            I => \N__52759\
        );

    \I__12767\ : InMux
    port map (
            O => \N__52819\,
            I => \N__52743\
        );

    \I__12766\ : LocalMux
    port map (
            O => \N__52806\,
            I => \N__52740\
        );

    \I__12765\ : Span4Mux_v
    port map (
            O => \N__52801\,
            I => \N__52735\
        );

    \I__12764\ : Span4Mux_h
    port map (
            O => \N__52796\,
            I => \N__52735\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__52793\,
            I => \N__52722\
        );

    \I__12762\ : LocalMux
    port map (
            O => \N__52788\,
            I => \N__52722\
        );

    \I__12761\ : LocalMux
    port map (
            O => \N__52779\,
            I => \N__52722\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__52774\,
            I => \N__52722\
        );

    \I__12759\ : Span4Mux_h
    port map (
            O => \N__52769\,
            I => \N__52722\
        );

    \I__12758\ : Span4Mux_v
    port map (
            O => \N__52764\,
            I => \N__52722\
        );

    \I__12757\ : Span4Mux_v
    port map (
            O => \N__52759\,
            I => \N__52717\
        );

    \I__12756\ : InMux
    port map (
            O => \N__52758\,
            I => \N__52710\
        );

    \I__12755\ : InMux
    port map (
            O => \N__52757\,
            I => \N__52710\
        );

    \I__12754\ : InMux
    port map (
            O => \N__52756\,
            I => \N__52710\
        );

    \I__12753\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52703\
        );

    \I__12752\ : InMux
    port map (
            O => \N__52754\,
            I => \N__52696\
        );

    \I__12751\ : InMux
    port map (
            O => \N__52753\,
            I => \N__52696\
        );

    \I__12750\ : InMux
    port map (
            O => \N__52752\,
            I => \N__52696\
        );

    \I__12749\ : InMux
    port map (
            O => \N__52751\,
            I => \N__52683\
        );

    \I__12748\ : InMux
    port map (
            O => \N__52750\,
            I => \N__52683\
        );

    \I__12747\ : InMux
    port map (
            O => \N__52749\,
            I => \N__52683\
        );

    \I__12746\ : InMux
    port map (
            O => \N__52748\,
            I => \N__52683\
        );

    \I__12745\ : InMux
    port map (
            O => \N__52747\,
            I => \N__52683\
        );

    \I__12744\ : InMux
    port map (
            O => \N__52746\,
            I => \N__52683\
        );

    \I__12743\ : LocalMux
    port map (
            O => \N__52743\,
            I => \N__52680\
        );

    \I__12742\ : Span4Mux_v
    port map (
            O => \N__52740\,
            I => \N__52675\
        );

    \I__12741\ : Span4Mux_h
    port map (
            O => \N__52735\,
            I => \N__52675\
        );

    \I__12740\ : Span4Mux_h
    port map (
            O => \N__52722\,
            I => \N__52672\
        );

    \I__12739\ : InMux
    port map (
            O => \N__52721\,
            I => \N__52667\
        );

    \I__12738\ : InMux
    port map (
            O => \N__52720\,
            I => \N__52667\
        );

    \I__12737\ : Span4Mux_h
    port map (
            O => \N__52717\,
            I => \N__52662\
        );

    \I__12736\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52662\
        );

    \I__12735\ : InMux
    port map (
            O => \N__52709\,
            I => \N__52653\
        );

    \I__12734\ : InMux
    port map (
            O => \N__52708\,
            I => \N__52653\
        );

    \I__12733\ : InMux
    port map (
            O => \N__52707\,
            I => \N__52653\
        );

    \I__12732\ : InMux
    port map (
            O => \N__52706\,
            I => \N__52653\
        );

    \I__12731\ : LocalMux
    port map (
            O => \N__52703\,
            I => adc_state_0_adj_1418
        );

    \I__12730\ : LocalMux
    port map (
            O => \N__52696\,
            I => adc_state_0_adj_1418
        );

    \I__12729\ : LocalMux
    port map (
            O => \N__52683\,
            I => adc_state_0_adj_1418
        );

    \I__12728\ : Odrv4
    port map (
            O => \N__52680\,
            I => adc_state_0_adj_1418
        );

    \I__12727\ : Odrv4
    port map (
            O => \N__52675\,
            I => adc_state_0_adj_1418
        );

    \I__12726\ : Odrv4
    port map (
            O => \N__52672\,
            I => adc_state_0_adj_1418
        );

    \I__12725\ : LocalMux
    port map (
            O => \N__52667\,
            I => adc_state_0_adj_1418
        );

    \I__12724\ : Odrv4
    port map (
            O => \N__52662\,
            I => adc_state_0_adj_1418
        );

    \I__12723\ : LocalMux
    port map (
            O => \N__52653\,
            I => adc_state_0_adj_1418
        );

    \I__12722\ : CascadeMux
    port map (
            O => \N__52634\,
            I => \N__52630\
        );

    \I__12721\ : CascadeMux
    port map (
            O => \N__52633\,
            I => \N__52627\
        );

    \I__12720\ : InMux
    port map (
            O => \N__52630\,
            I => \N__52623\
        );

    \I__12719\ : InMux
    port map (
            O => \N__52627\,
            I => \N__52618\
        );

    \I__12718\ : InMux
    port map (
            O => \N__52626\,
            I => \N__52618\
        );

    \I__12717\ : LocalMux
    port map (
            O => \N__52623\,
            I => cmd_rdadctmp_17_adj_1433
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__52618\,
            I => cmd_rdadctmp_17_adj_1433
        );

    \I__12715\ : InMux
    port map (
            O => \N__52613\,
            I => \N__52610\
        );

    \I__12714\ : LocalMux
    port map (
            O => \N__52610\,
            I => \N__52606\
        );

    \I__12713\ : InMux
    port map (
            O => \N__52609\,
            I => \N__52603\
        );

    \I__12712\ : Span4Mux_h
    port map (
            O => \N__52606\,
            I => \N__52599\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52596\
        );

    \I__12710\ : InMux
    port map (
            O => \N__52602\,
            I => \N__52593\
        );

    \I__12709\ : Span4Mux_v
    port map (
            O => \N__52599\,
            I => \N__52588\
        );

    \I__12708\ : Span4Mux_h
    port map (
            O => \N__52596\,
            I => \N__52588\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__52593\,
            I => buf_adcdata_iac_9
        );

    \I__12706\ : Odrv4
    port map (
            O => \N__52588\,
            I => buf_adcdata_iac_9
        );

    \I__12705\ : InMux
    port map (
            O => \N__52583\,
            I => \N__52580\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__52580\,
            I => \N__52577\
        );

    \I__12703\ : Span4Mux_h
    port map (
            O => \N__52577\,
            I => \N__52574\
        );

    \I__12702\ : Odrv4
    port map (
            O => \N__52574\,
            I => buf_data_iac_12
        );

    \I__12701\ : CascadeMux
    port map (
            O => \N__52571\,
            I => \N__52568\
        );

    \I__12700\ : InMux
    port map (
            O => \N__52568\,
            I => \N__52565\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__52565\,
            I => \N__52562\
        );

    \I__12698\ : Span4Mux_h
    port map (
            O => \N__52562\,
            I => \N__52559\
        );

    \I__12697\ : Span4Mux_h
    port map (
            O => \N__52559\,
            I => \N__52556\
        );

    \I__12696\ : Odrv4
    port map (
            O => \N__52556\,
            I => n21230
        );

    \I__12695\ : InMux
    port map (
            O => \N__52553\,
            I => \N__52550\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__52550\,
            I => \N__52547\
        );

    \I__12693\ : Span4Mux_h
    port map (
            O => \N__52547\,
            I => \N__52544\
        );

    \I__12692\ : Odrv4
    port map (
            O => \N__52544\,
            I => buf_data_iac_13
        );

    \I__12691\ : InMux
    port map (
            O => \N__52541\,
            I => \N__52538\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__52538\,
            I => \N__52535\
        );

    \I__12689\ : Span4Mux_v
    port map (
            O => \N__52535\,
            I => \N__52532\
        );

    \I__12688\ : Span4Mux_h
    port map (
            O => \N__52532\,
            I => \N__52529\
        );

    \I__12687\ : Odrv4
    port map (
            O => \N__52529\,
            I => n21297
        );

    \I__12686\ : SRMux
    port map (
            O => \N__52526\,
            I => \N__52523\
        );

    \I__12685\ : LocalMux
    port map (
            O => \N__52523\,
            I => \N__52520\
        );

    \I__12684\ : Span4Mux_h
    port map (
            O => \N__52520\,
            I => \N__52517\
        );

    \I__12683\ : Span4Mux_v
    port map (
            O => \N__52517\,
            I => \N__52514\
        );

    \I__12682\ : Odrv4
    port map (
            O => \N__52514\,
            I => \comm_spi.DOUT_7__N_747\
        );

    \I__12681\ : CascadeMux
    port map (
            O => \N__52511\,
            I => \N__52508\
        );

    \I__12680\ : InMux
    port map (
            O => \N__52508\,
            I => \N__52500\
        );

    \I__12679\ : InMux
    port map (
            O => \N__52507\,
            I => \N__52500\
        );

    \I__12678\ : CascadeMux
    port map (
            O => \N__52506\,
            I => \N__52497\
        );

    \I__12677\ : InMux
    port map (
            O => \N__52505\,
            I => \N__52494\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__52500\,
            I => \N__52490\
        );

    \I__12675\ : InMux
    port map (
            O => \N__52497\,
            I => \N__52486\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__52494\,
            I => \N__52483\
        );

    \I__12673\ : InMux
    port map (
            O => \N__52493\,
            I => \N__52480\
        );

    \I__12672\ : Span4Mux_v
    port map (
            O => \N__52490\,
            I => \N__52477\
        );

    \I__12671\ : InMux
    port map (
            O => \N__52489\,
            I => \N__52474\
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__52486\,
            I => \N__52471\
        );

    \I__12669\ : Span4Mux_v
    port map (
            O => \N__52483\,
            I => \N__52468\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__52480\,
            I => \N__52465\
        );

    \I__12667\ : Span4Mux_h
    port map (
            O => \N__52477\,
            I => \N__52460\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__52474\,
            I => \N__52460\
        );

    \I__12665\ : Span4Mux_v
    port map (
            O => \N__52471\,
            I => \N__52457\
        );

    \I__12664\ : Sp12to4
    port map (
            O => \N__52468\,
            I => \N__52454\
        );

    \I__12663\ : Span4Mux_v
    port map (
            O => \N__52465\,
            I => \N__52451\
        );

    \I__12662\ : Span4Mux_v
    port map (
            O => \N__52460\,
            I => \N__52448\
        );

    \I__12661\ : Odrv4
    port map (
            O => \N__52457\,
            I => comm_buf_1_6
        );

    \I__12660\ : Odrv12
    port map (
            O => \N__52454\,
            I => comm_buf_1_6
        );

    \I__12659\ : Odrv4
    port map (
            O => \N__52451\,
            I => comm_buf_1_6
        );

    \I__12658\ : Odrv4
    port map (
            O => \N__52448\,
            I => comm_buf_1_6
        );

    \I__12657\ : InMux
    port map (
            O => \N__52439\,
            I => \N__52421\
        );

    \I__12656\ : InMux
    port map (
            O => \N__52438\,
            I => \N__52421\
        );

    \I__12655\ : InMux
    port map (
            O => \N__52437\,
            I => \N__52421\
        );

    \I__12654\ : InMux
    port map (
            O => \N__52436\,
            I => \N__52421\
        );

    \I__12653\ : InMux
    port map (
            O => \N__52435\,
            I => \N__52421\
        );

    \I__12652\ : InMux
    port map (
            O => \N__52434\,
            I => \N__52417\
        );

    \I__12651\ : InMux
    port map (
            O => \N__52433\,
            I => \N__52413\
        );

    \I__12650\ : InMux
    port map (
            O => \N__52432\,
            I => \N__52403\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__52421\,
            I => \N__52400\
        );

    \I__12648\ : InMux
    port map (
            O => \N__52420\,
            I => \N__52397\
        );

    \I__12647\ : LocalMux
    port map (
            O => \N__52417\,
            I => \N__52394\
        );

    \I__12646\ : InMux
    port map (
            O => \N__52416\,
            I => \N__52384\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__52413\,
            I => \N__52381\
        );

    \I__12644\ : InMux
    port map (
            O => \N__52412\,
            I => \N__52371\
        );

    \I__12643\ : InMux
    port map (
            O => \N__52411\,
            I => \N__52371\
        );

    \I__12642\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52361\
        );

    \I__12641\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52356\
        );

    \I__12640\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52356\
        );

    \I__12639\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52353\
        );

    \I__12638\ : CascadeMux
    port map (
            O => \N__52406\,
            I => \N__52350\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__52403\,
            I => \N__52345\
        );

    \I__12636\ : Span4Mux_v
    port map (
            O => \N__52400\,
            I => \N__52342\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__52397\,
            I => \N__52339\
        );

    \I__12634\ : Span4Mux_h
    port map (
            O => \N__52394\,
            I => \N__52336\
        );

    \I__12633\ : InMux
    port map (
            O => \N__52393\,
            I => \N__52327\
        );

    \I__12632\ : InMux
    port map (
            O => \N__52392\,
            I => \N__52327\
        );

    \I__12631\ : InMux
    port map (
            O => \N__52391\,
            I => \N__52327\
        );

    \I__12630\ : InMux
    port map (
            O => \N__52390\,
            I => \N__52327\
        );

    \I__12629\ : InMux
    port map (
            O => \N__52389\,
            I => \N__52319\
        );

    \I__12628\ : InMux
    port map (
            O => \N__52388\,
            I => \N__52319\
        );

    \I__12627\ : InMux
    port map (
            O => \N__52387\,
            I => \N__52319\
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__52384\,
            I => \N__52314\
        );

    \I__12625\ : Span4Mux_h
    port map (
            O => \N__52381\,
            I => \N__52314\
        );

    \I__12624\ : InMux
    port map (
            O => \N__52380\,
            I => \N__52307\
        );

    \I__12623\ : InMux
    port map (
            O => \N__52379\,
            I => \N__52307\
        );

    \I__12622\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52307\
        );

    \I__12621\ : InMux
    port map (
            O => \N__52377\,
            I => \N__52297\
        );

    \I__12620\ : InMux
    port map (
            O => \N__52376\,
            I => \N__52297\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__52371\,
            I => \N__52294\
        );

    \I__12618\ : InMux
    port map (
            O => \N__52370\,
            I => \N__52289\
        );

    \I__12617\ : InMux
    port map (
            O => \N__52369\,
            I => \N__52289\
        );

    \I__12616\ : InMux
    port map (
            O => \N__52368\,
            I => \N__52286\
        );

    \I__12615\ : InMux
    port map (
            O => \N__52367\,
            I => \N__52283\
        );

    \I__12614\ : InMux
    port map (
            O => \N__52366\,
            I => \N__52280\
        );

    \I__12613\ : InMux
    port map (
            O => \N__52365\,
            I => \N__52275\
        );

    \I__12612\ : InMux
    port map (
            O => \N__52364\,
            I => \N__52275\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__52361\,
            I => \N__52270\
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__52356\,
            I => \N__52270\
        );

    \I__12609\ : LocalMux
    port map (
            O => \N__52353\,
            I => \N__52267\
        );

    \I__12608\ : InMux
    port map (
            O => \N__52350\,
            I => \N__52260\
        );

    \I__12607\ : InMux
    port map (
            O => \N__52349\,
            I => \N__52260\
        );

    \I__12606\ : InMux
    port map (
            O => \N__52348\,
            I => \N__52260\
        );

    \I__12605\ : Span4Mux_v
    port map (
            O => \N__52345\,
            I => \N__52254\
        );

    \I__12604\ : Span4Mux_h
    port map (
            O => \N__52342\,
            I => \N__52254\
        );

    \I__12603\ : Span4Mux_h
    port map (
            O => \N__52339\,
            I => \N__52247\
        );

    \I__12602\ : Span4Mux_v
    port map (
            O => \N__52336\,
            I => \N__52247\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__52327\,
            I => \N__52247\
        );

    \I__12600\ : InMux
    port map (
            O => \N__52326\,
            I => \N__52244\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__52319\,
            I => \N__52237\
        );

    \I__12598\ : Sp12to4
    port map (
            O => \N__52314\,
            I => \N__52237\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__52307\,
            I => \N__52237\
        );

    \I__12596\ : InMux
    port map (
            O => \N__52306\,
            I => \N__52232\
        );

    \I__12595\ : InMux
    port map (
            O => \N__52305\,
            I => \N__52232\
        );

    \I__12594\ : InMux
    port map (
            O => \N__52304\,
            I => \N__52225\
        );

    \I__12593\ : InMux
    port map (
            O => \N__52303\,
            I => \N__52225\
        );

    \I__12592\ : InMux
    port map (
            O => \N__52302\,
            I => \N__52225\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__52297\,
            I => \N__52216\
        );

    \I__12590\ : Span4Mux_v
    port map (
            O => \N__52294\,
            I => \N__52216\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__52289\,
            I => \N__52216\
        );

    \I__12588\ : LocalMux
    port map (
            O => \N__52286\,
            I => \N__52216\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__52283\,
            I => \N__52203\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__52280\,
            I => \N__52203\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__52275\,
            I => \N__52203\
        );

    \I__12584\ : Sp12to4
    port map (
            O => \N__52270\,
            I => \N__52203\
        );

    \I__12583\ : Span12Mux_h
    port map (
            O => \N__52267\,
            I => \N__52203\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__52260\,
            I => \N__52203\
        );

    \I__12581\ : InMux
    port map (
            O => \N__52259\,
            I => \N__52200\
        );

    \I__12580\ : Span4Mux_h
    port map (
            O => \N__52254\,
            I => \N__52195\
        );

    \I__12579\ : Span4Mux_v
    port map (
            O => \N__52247\,
            I => \N__52195\
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__52244\,
            I => \N__52190\
        );

    \I__12577\ : Span12Mux_v
    port map (
            O => \N__52237\,
            I => \N__52190\
        );

    \I__12576\ : LocalMux
    port map (
            O => \N__52232\,
            I => comm_state_2
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__52225\,
            I => comm_state_2
        );

    \I__12574\ : Odrv4
    port map (
            O => \N__52216\,
            I => comm_state_2
        );

    \I__12573\ : Odrv12
    port map (
            O => \N__52203\,
            I => comm_state_2
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__52200\,
            I => comm_state_2
        );

    \I__12571\ : Odrv4
    port map (
            O => \N__52195\,
            I => comm_state_2
        );

    \I__12570\ : Odrv12
    port map (
            O => \N__52190\,
            I => comm_state_2
        );

    \I__12569\ : InMux
    port map (
            O => \N__52175\,
            I => \N__52171\
        );

    \I__12568\ : InMux
    port map (
            O => \N__52174\,
            I => \N__52168\
        );

    \I__12567\ : LocalMux
    port map (
            O => \N__52171\,
            I => \N__52165\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__52168\,
            I => \N__52160\
        );

    \I__12565\ : Span4Mux_h
    port map (
            O => \N__52165\,
            I => \N__52160\
        );

    \I__12564\ : Odrv4
    port map (
            O => \N__52160\,
            I => n14_adj_1547
        );

    \I__12563\ : CascadeMux
    port map (
            O => \N__52157\,
            I => \N__52154\
        );

    \I__12562\ : InMux
    port map (
            O => \N__52154\,
            I => \N__52150\
        );

    \I__12561\ : InMux
    port map (
            O => \N__52153\,
            I => \N__52147\
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__52150\,
            I => \N__52144\
        );

    \I__12559\ : LocalMux
    port map (
            O => \N__52147\,
            I => \N__52140\
        );

    \I__12558\ : Span4Mux_v
    port map (
            O => \N__52144\,
            I => \N__52137\
        );

    \I__12557\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52134\
        );

    \I__12556\ : Span12Mux_s10_h
    port map (
            O => \N__52140\,
            I => \N__52131\
        );

    \I__12555\ : Span4Mux_h
    port map (
            O => \N__52137\,
            I => \N__52128\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__52134\,
            I => buf_adcdata_iac_8
        );

    \I__12553\ : Odrv12
    port map (
            O => \N__52131\,
            I => buf_adcdata_iac_8
        );

    \I__12552\ : Odrv4
    port map (
            O => \N__52128\,
            I => buf_adcdata_iac_8
        );

    \I__12551\ : CascadeMux
    port map (
            O => \N__52121\,
            I => \N__52117\
        );

    \I__12550\ : CascadeMux
    port map (
            O => \N__52120\,
            I => \N__52114\
        );

    \I__12549\ : InMux
    port map (
            O => \N__52117\,
            I => \N__52109\
        );

    \I__12548\ : InMux
    port map (
            O => \N__52114\,
            I => \N__52109\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__52109\,
            I => \N__52106\
        );

    \I__12546\ : Span12Mux_v
    port map (
            O => \N__52106\,
            I => \N__52102\
        );

    \I__12545\ : InMux
    port map (
            O => \N__52105\,
            I => \N__52099\
        );

    \I__12544\ : Odrv12
    port map (
            O => \N__52102\,
            I => cmd_rdadctmp_16_adj_1434
        );

    \I__12543\ : LocalMux
    port map (
            O => \N__52099\,
            I => cmd_rdadctmp_16_adj_1434
        );

    \I__12542\ : InMux
    port map (
            O => \N__52094\,
            I => \N__52091\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__52091\,
            I => \N__52082\
        );

    \I__12540\ : InMux
    port map (
            O => \N__52090\,
            I => \N__52079\
        );

    \I__12539\ : InMux
    port map (
            O => \N__52089\,
            I => \N__52068\
        );

    \I__12538\ : InMux
    port map (
            O => \N__52088\,
            I => \N__52065\
        );

    \I__12537\ : InMux
    port map (
            O => \N__52087\,
            I => \N__52058\
        );

    \I__12536\ : InMux
    port map (
            O => \N__52086\,
            I => \N__52058\
        );

    \I__12535\ : InMux
    port map (
            O => \N__52085\,
            I => \N__52058\
        );

    \I__12534\ : Span4Mux_h
    port map (
            O => \N__52082\,
            I => \N__52053\
        );

    \I__12533\ : LocalMux
    port map (
            O => \N__52079\,
            I => \N__52053\
        );

    \I__12532\ : InMux
    port map (
            O => \N__52078\,
            I => \N__52048\
        );

    \I__12531\ : InMux
    port map (
            O => \N__52077\,
            I => \N__52048\
        );

    \I__12530\ : InMux
    port map (
            O => \N__52076\,
            I => \N__52043\
        );

    \I__12529\ : InMux
    port map (
            O => \N__52075\,
            I => \N__52040\
        );

    \I__12528\ : InMux
    port map (
            O => \N__52074\,
            I => \N__52031\
        );

    \I__12527\ : InMux
    port map (
            O => \N__52073\,
            I => \N__52031\
        );

    \I__12526\ : InMux
    port map (
            O => \N__52072\,
            I => \N__52031\
        );

    \I__12525\ : InMux
    port map (
            O => \N__52071\,
            I => \N__52031\
        );

    \I__12524\ : LocalMux
    port map (
            O => \N__52068\,
            I => \N__52028\
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__52065\,
            I => \N__52023\
        );

    \I__12522\ : LocalMux
    port map (
            O => \N__52058\,
            I => \N__52023\
        );

    \I__12521\ : Span4Mux_v
    port map (
            O => \N__52053\,
            I => \N__52020\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__52048\,
            I => \N__52017\
        );

    \I__12519\ : InMux
    port map (
            O => \N__52047\,
            I => \N__52009\
        );

    \I__12518\ : InMux
    port map (
            O => \N__52046\,
            I => \N__52009\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__52043\,
            I => \N__52006\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__52040\,
            I => \N__51999\
        );

    \I__12515\ : LocalMux
    port map (
            O => \N__52031\,
            I => \N__51994\
        );

    \I__12514\ : Sp12to4
    port map (
            O => \N__52028\,
            I => \N__51994\
        );

    \I__12513\ : Span4Mux_v
    port map (
            O => \N__52023\,
            I => \N__51991\
        );

    \I__12512\ : Span4Mux_h
    port map (
            O => \N__52020\,
            I => \N__51988\
        );

    \I__12511\ : Span4Mux_v
    port map (
            O => \N__52017\,
            I => \N__51985\
        );

    \I__12510\ : InMux
    port map (
            O => \N__52016\,
            I => \N__51974\
        );

    \I__12509\ : InMux
    port map (
            O => \N__52015\,
            I => \N__51969\
        );

    \I__12508\ : InMux
    port map (
            O => \N__52014\,
            I => \N__51969\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__52009\,
            I => \N__51964\
        );

    \I__12506\ : Span4Mux_h
    port map (
            O => \N__52006\,
            I => \N__51964\
        );

    \I__12505\ : InMux
    port map (
            O => \N__52005\,
            I => \N__51959\
        );

    \I__12504\ : InMux
    port map (
            O => \N__52004\,
            I => \N__51959\
        );

    \I__12503\ : InMux
    port map (
            O => \N__52003\,
            I => \N__51954\
        );

    \I__12502\ : InMux
    port map (
            O => \N__52002\,
            I => \N__51954\
        );

    \I__12501\ : Sp12to4
    port map (
            O => \N__51999\,
            I => \N__51947\
        );

    \I__12500\ : Span12Mux_v
    port map (
            O => \N__51994\,
            I => \N__51947\
        );

    \I__12499\ : Sp12to4
    port map (
            O => \N__51991\,
            I => \N__51947\
        );

    \I__12498\ : Sp12to4
    port map (
            O => \N__51988\,
            I => \N__51942\
        );

    \I__12497\ : Sp12to4
    port map (
            O => \N__51985\,
            I => \N__51942\
        );

    \I__12496\ : InMux
    port map (
            O => \N__51984\,
            I => \N__51937\
        );

    \I__12495\ : InMux
    port map (
            O => \N__51983\,
            I => \N__51937\
        );

    \I__12494\ : InMux
    port map (
            O => \N__51982\,
            I => \N__51932\
        );

    \I__12493\ : InMux
    port map (
            O => \N__51981\,
            I => \N__51932\
        );

    \I__12492\ : InMux
    port map (
            O => \N__51980\,
            I => \N__51923\
        );

    \I__12491\ : InMux
    port map (
            O => \N__51979\,
            I => \N__51923\
        );

    \I__12490\ : InMux
    port map (
            O => \N__51978\,
            I => \N__51923\
        );

    \I__12489\ : InMux
    port map (
            O => \N__51977\,
            I => \N__51923\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__51974\,
            I => \N__51920\
        );

    \I__12487\ : LocalMux
    port map (
            O => \N__51969\,
            I => \N__51915\
        );

    \I__12486\ : Span4Mux_h
    port map (
            O => \N__51964\,
            I => \N__51915\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__51959\,
            I => \N__51908\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__51954\,
            I => \N__51908\
        );

    \I__12483\ : Span12Mux_h
    port map (
            O => \N__51947\,
            I => \N__51908\
        );

    \I__12482\ : Span12Mux_h
    port map (
            O => \N__51942\,
            I => \N__51905\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__51937\,
            I => n12663
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__51932\,
            I => n12663
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__51923\,
            I => n12663
        );

    \I__12478\ : Odrv4
    port map (
            O => \N__51920\,
            I => n12663
        );

    \I__12477\ : Odrv4
    port map (
            O => \N__51915\,
            I => n12663
        );

    \I__12476\ : Odrv12
    port map (
            O => \N__51908\,
            I => n12663
        );

    \I__12475\ : Odrv12
    port map (
            O => \N__51905\,
            I => n12663
        );

    \I__12474\ : CascadeMux
    port map (
            O => \N__51890\,
            I => \N__51886\
        );

    \I__12473\ : InMux
    port map (
            O => \N__51889\,
            I => \N__51878\
        );

    \I__12472\ : InMux
    port map (
            O => \N__51886\,
            I => \N__51878\
        );

    \I__12471\ : InMux
    port map (
            O => \N__51885\,
            I => \N__51878\
        );

    \I__12470\ : LocalMux
    port map (
            O => \N__51878\,
            I => cmd_rdadctmp_18_adj_1432
        );

    \I__12469\ : InMux
    port map (
            O => \N__51875\,
            I => \N__51870\
        );

    \I__12468\ : CascadeMux
    port map (
            O => \N__51874\,
            I => \N__51867\
        );

    \I__12467\ : CascadeMux
    port map (
            O => \N__51873\,
            I => \N__51864\
        );

    \I__12466\ : LocalMux
    port map (
            O => \N__51870\,
            I => \N__51861\
        );

    \I__12465\ : InMux
    port map (
            O => \N__51867\,
            I => \N__51858\
        );

    \I__12464\ : InMux
    port map (
            O => \N__51864\,
            I => \N__51855\
        );

    \I__12463\ : Span12Mux_v
    port map (
            O => \N__51861\,
            I => \N__51852\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__51858\,
            I => buf_adcdata_iac_10
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__51855\,
            I => buf_adcdata_iac_10
        );

    \I__12460\ : Odrv12
    port map (
            O => \N__51852\,
            I => buf_adcdata_iac_10
        );

    \I__12459\ : CascadeMux
    port map (
            O => \N__51845\,
            I => \N__51835\
        );

    \I__12458\ : CascadeMux
    port map (
            O => \N__51844\,
            I => \N__51832\
        );

    \I__12457\ : CascadeMux
    port map (
            O => \N__51843\,
            I => \N__51829\
        );

    \I__12456\ : InMux
    port map (
            O => \N__51842\,
            I => \N__51820\
        );

    \I__12455\ : InMux
    port map (
            O => \N__51841\,
            I => \N__51820\
        );

    \I__12454\ : InMux
    port map (
            O => \N__51840\,
            I => \N__51817\
        );

    \I__12453\ : InMux
    port map (
            O => \N__51839\,
            I => \N__51814\
        );

    \I__12452\ : CascadeMux
    port map (
            O => \N__51838\,
            I => \N__51811\
        );

    \I__12451\ : InMux
    port map (
            O => \N__51835\,
            I => \N__51804\
        );

    \I__12450\ : InMux
    port map (
            O => \N__51832\,
            I => \N__51804\
        );

    \I__12449\ : InMux
    port map (
            O => \N__51829\,
            I => \N__51804\
        );

    \I__12448\ : InMux
    port map (
            O => \N__51828\,
            I => \N__51801\
        );

    \I__12447\ : InMux
    port map (
            O => \N__51827\,
            I => \N__51794\
        );

    \I__12446\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51794\
        );

    \I__12445\ : InMux
    port map (
            O => \N__51825\,
            I => \N__51794\
        );

    \I__12444\ : LocalMux
    port map (
            O => \N__51820\,
            I => \N__51789\
        );

    \I__12443\ : LocalMux
    port map (
            O => \N__51817\,
            I => \N__51789\
        );

    \I__12442\ : LocalMux
    port map (
            O => \N__51814\,
            I => \N__51786\
        );

    \I__12441\ : InMux
    port map (
            O => \N__51811\,
            I => \N__51783\
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__51804\,
            I => \N__51777\
        );

    \I__12439\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51777\
        );

    \I__12438\ : LocalMux
    port map (
            O => \N__51794\,
            I => \N__51774\
        );

    \I__12437\ : Span4Mux_v
    port map (
            O => \N__51789\,
            I => \N__51767\
        );

    \I__12436\ : Span4Mux_h
    port map (
            O => \N__51786\,
            I => \N__51767\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__51783\,
            I => \N__51767\
        );

    \I__12434\ : CascadeMux
    port map (
            O => \N__51782\,
            I => \N__51763\
        );

    \I__12433\ : Span4Mux_v
    port map (
            O => \N__51777\,
            I => \N__51759\
        );

    \I__12432\ : Span4Mux_v
    port map (
            O => \N__51774\,
            I => \N__51756\
        );

    \I__12431\ : Span4Mux_v
    port map (
            O => \N__51767\,
            I => \N__51753\
        );

    \I__12430\ : InMux
    port map (
            O => \N__51766\,
            I => \N__51748\
        );

    \I__12429\ : InMux
    port map (
            O => \N__51763\,
            I => \N__51748\
        );

    \I__12428\ : CascadeMux
    port map (
            O => \N__51762\,
            I => \N__51742\
        );

    \I__12427\ : Sp12to4
    port map (
            O => \N__51759\,
            I => \N__51738\
        );

    \I__12426\ : Sp12to4
    port map (
            O => \N__51756\,
            I => \N__51735\
        );

    \I__12425\ : Span4Mux_h
    port map (
            O => \N__51753\,
            I => \N__51732\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__51748\,
            I => \N__51729\
        );

    \I__12423\ : InMux
    port map (
            O => \N__51747\,
            I => \N__51724\
        );

    \I__12422\ : InMux
    port map (
            O => \N__51746\,
            I => \N__51724\
        );

    \I__12421\ : InMux
    port map (
            O => \N__51745\,
            I => \N__51717\
        );

    \I__12420\ : InMux
    port map (
            O => \N__51742\,
            I => \N__51717\
        );

    \I__12419\ : InMux
    port map (
            O => \N__51741\,
            I => \N__51717\
        );

    \I__12418\ : Span12Mux_h
    port map (
            O => \N__51738\,
            I => \N__51714\
        );

    \I__12417\ : Span12Mux_s10_h
    port map (
            O => \N__51735\,
            I => \N__51703\
        );

    \I__12416\ : Sp12to4
    port map (
            O => \N__51732\,
            I => \N__51703\
        );

    \I__12415\ : Sp12to4
    port map (
            O => \N__51729\,
            I => \N__51703\
        );

    \I__12414\ : LocalMux
    port map (
            O => \N__51724\,
            I => \N__51703\
        );

    \I__12413\ : LocalMux
    port map (
            O => \N__51717\,
            I => \N__51703\
        );

    \I__12412\ : Span12Mux_v
    port map (
            O => \N__51714\,
            I => \N__51700\
        );

    \I__12411\ : Span12Mux_v
    port map (
            O => \N__51703\,
            I => \N__51697\
        );

    \I__12410\ : Odrv12
    port map (
            O => \N__51700\,
            I => \ICE_SPI_CE0\
        );

    \I__12409\ : Odrv12
    port map (
            O => \N__51697\,
            I => \ICE_SPI_CE0\
        );

    \I__12408\ : InMux
    port map (
            O => \N__51692\,
            I => \N__51683\
        );

    \I__12407\ : InMux
    port map (
            O => \N__51691\,
            I => \N__51683\
        );

    \I__12406\ : InMux
    port map (
            O => \N__51690\,
            I => \N__51680\
        );

    \I__12405\ : InMux
    port map (
            O => \N__51689\,
            I => \N__51677\
        );

    \I__12404\ : InMux
    port map (
            O => \N__51688\,
            I => \N__51674\
        );

    \I__12403\ : LocalMux
    port map (
            O => \N__51683\,
            I => \N__51666\
        );

    \I__12402\ : LocalMux
    port map (
            O => \N__51680\,
            I => \N__51663\
        );

    \I__12401\ : LocalMux
    port map (
            O => \N__51677\,
            I => \N__51658\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__51674\,
            I => \N__51658\
        );

    \I__12399\ : InMux
    port map (
            O => \N__51673\,
            I => \N__51653\
        );

    \I__12398\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51653\
        );

    \I__12397\ : InMux
    port map (
            O => \N__51671\,
            I => \N__51648\
        );

    \I__12396\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51648\
        );

    \I__12395\ : CascadeMux
    port map (
            O => \N__51669\,
            I => \N__51643\
        );

    \I__12394\ : Span4Mux_h
    port map (
            O => \N__51666\,
            I => \N__51639\
        );

    \I__12393\ : Span4Mux_v
    port map (
            O => \N__51663\,
            I => \N__51632\
        );

    \I__12392\ : Span4Mux_v
    port map (
            O => \N__51658\,
            I => \N__51632\
        );

    \I__12391\ : LocalMux
    port map (
            O => \N__51653\,
            I => \N__51632\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__51648\,
            I => \N__51629\
        );

    \I__12389\ : InMux
    port map (
            O => \N__51647\,
            I => \N__51620\
        );

    \I__12388\ : InMux
    port map (
            O => \N__51646\,
            I => \N__51620\
        );

    \I__12387\ : InMux
    port map (
            O => \N__51643\,
            I => \N__51620\
        );

    \I__12386\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51620\
        );

    \I__12385\ : Odrv4
    port map (
            O => \N__51639\,
            I => comm_data_vld
        );

    \I__12384\ : Odrv4
    port map (
            O => \N__51632\,
            I => comm_data_vld
        );

    \I__12383\ : Odrv4
    port map (
            O => \N__51629\,
            I => comm_data_vld
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__51620\,
            I => comm_data_vld
        );

    \I__12381\ : InMux
    port map (
            O => \N__51611\,
            I => \N__51608\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__51608\,
            I => n21129
        );

    \I__12379\ : CascadeMux
    port map (
            O => \N__51605\,
            I => \N__51602\
        );

    \I__12378\ : InMux
    port map (
            O => \N__51602\,
            I => \N__51599\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__51599\,
            I => \N__51596\
        );

    \I__12376\ : Odrv4
    port map (
            O => \N__51596\,
            I => n20740
        );

    \I__12375\ : CascadeMux
    port map (
            O => \N__51593\,
            I => \n11363_cascade_\
        );

    \I__12374\ : CascadeMux
    port map (
            O => \N__51590\,
            I => \N__51586\
        );

    \I__12373\ : InMux
    port map (
            O => \N__51589\,
            I => \N__51581\
        );

    \I__12372\ : InMux
    port map (
            O => \N__51586\,
            I => \N__51574\
        );

    \I__12371\ : InMux
    port map (
            O => \N__51585\,
            I => \N__51574\
        );

    \I__12370\ : InMux
    port map (
            O => \N__51584\,
            I => \N__51574\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__51581\,
            I => \N__51570\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__51574\,
            I => \N__51565\
        );

    \I__12367\ : CascadeMux
    port map (
            O => \N__51573\,
            I => \N__51562\
        );

    \I__12366\ : Span4Mux_v
    port map (
            O => \N__51570\,
            I => \N__51559\
        );

    \I__12365\ : CascadeMux
    port map (
            O => \N__51569\,
            I => \N__51556\
        );

    \I__12364\ : InMux
    port map (
            O => \N__51568\,
            I => \N__51553\
        );

    \I__12363\ : Span4Mux_h
    port map (
            O => \N__51565\,
            I => \N__51546\
        );

    \I__12362\ : InMux
    port map (
            O => \N__51562\,
            I => \N__51543\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__51559\,
            I => \N__51539\
        );

    \I__12360\ : InMux
    port map (
            O => \N__51556\,
            I => \N__51536\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__51553\,
            I => \N__51533\
        );

    \I__12358\ : InMux
    port map (
            O => \N__51552\,
            I => \N__51530\
        );

    \I__12357\ : InMux
    port map (
            O => \N__51551\,
            I => \N__51527\
        );

    \I__12356\ : InMux
    port map (
            O => \N__51550\,
            I => \N__51522\
        );

    \I__12355\ : InMux
    port map (
            O => \N__51549\,
            I => \N__51522\
        );

    \I__12354\ : Span4Mux_h
    port map (
            O => \N__51546\,
            I => \N__51519\
        );

    \I__12353\ : LocalMux
    port map (
            O => \N__51543\,
            I => \N__51516\
        );

    \I__12352\ : InMux
    port map (
            O => \N__51542\,
            I => \N__51513\
        );

    \I__12351\ : Sp12to4
    port map (
            O => \N__51539\,
            I => \N__51508\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__51536\,
            I => \N__51508\
        );

    \I__12349\ : Span4Mux_h
    port map (
            O => \N__51533\,
            I => \N__51505\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__51530\,
            I => \N__51498\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__51527\,
            I => \N__51498\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__51522\,
            I => \N__51498\
        );

    \I__12345\ : Span4Mux_v
    port map (
            O => \N__51519\,
            I => \N__51493\
        );

    \I__12344\ : Span4Mux_h
    port map (
            O => \N__51516\,
            I => \N__51493\
        );

    \I__12343\ : LocalMux
    port map (
            O => \N__51513\,
            I => n12242
        );

    \I__12342\ : Odrv12
    port map (
            O => \N__51508\,
            I => n12242
        );

    \I__12341\ : Odrv4
    port map (
            O => \N__51505\,
            I => n12242
        );

    \I__12340\ : Odrv4
    port map (
            O => \N__51498\,
            I => n12242
        );

    \I__12339\ : Odrv4
    port map (
            O => \N__51493\,
            I => n12242
        );

    \I__12338\ : InMux
    port map (
            O => \N__51482\,
            I => \N__51478\
        );

    \I__12337\ : CascadeMux
    port map (
            O => \N__51481\,
            I => \N__51473\
        );

    \I__12336\ : LocalMux
    port map (
            O => \N__51478\,
            I => \N__51470\
        );

    \I__12335\ : InMux
    port map (
            O => \N__51477\,
            I => \N__51465\
        );

    \I__12334\ : InMux
    port map (
            O => \N__51476\,
            I => \N__51465\
        );

    \I__12333\ : InMux
    port map (
            O => \N__51473\,
            I => \N__51462\
        );

    \I__12332\ : Odrv4
    port map (
            O => \N__51470\,
            I => n12235
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__51465\,
            I => n12235
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__51462\,
            I => n12235
        );

    \I__12329\ : InMux
    port map (
            O => \N__51455\,
            I => \N__51452\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__51452\,
            I => \N__51449\
        );

    \I__12327\ : Span4Mux_h
    port map (
            O => \N__51449\,
            I => \N__51446\
        );

    \I__12326\ : Odrv4
    port map (
            O => \N__51446\,
            I => n11869
        );

    \I__12325\ : CEMux
    port map (
            O => \N__51443\,
            I => \N__51439\
        );

    \I__12324\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51436\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__51439\,
            I => \N__51432\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__51436\,
            I => \N__51429\
        );

    \I__12321\ : InMux
    port map (
            O => \N__51435\,
            I => \N__51426\
        );

    \I__12320\ : Span4Mux_h
    port map (
            O => \N__51432\,
            I => \N__51423\
        );

    \I__12319\ : Span4Mux_h
    port map (
            O => \N__51429\,
            I => \N__51418\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__51426\,
            I => \N__51418\
        );

    \I__12317\ : Span4Mux_v
    port map (
            O => \N__51423\,
            I => \N__51415\
        );

    \I__12316\ : Span4Mux_v
    port map (
            O => \N__51418\,
            I => \N__51412\
        );

    \I__12315\ : Odrv4
    port map (
            O => \N__51415\,
            I => n11876
        );

    \I__12314\ : Odrv4
    port map (
            O => \N__51412\,
            I => n11876
        );

    \I__12313\ : CascadeMux
    port map (
            O => \N__51407\,
            I => \N__51402\
        );

    \I__12312\ : InMux
    port map (
            O => \N__51406\,
            I => \N__51399\
        );

    \I__12311\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51395\
        );

    \I__12310\ : InMux
    port map (
            O => \N__51402\,
            I => \N__51390\
        );

    \I__12309\ : LocalMux
    port map (
            O => \N__51399\,
            I => \N__51387\
        );

    \I__12308\ : CascadeMux
    port map (
            O => \N__51398\,
            I => \N__51384\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__51395\,
            I => \N__51380\
        );

    \I__12306\ : InMux
    port map (
            O => \N__51394\,
            I => \N__51377\
        );

    \I__12305\ : InMux
    port map (
            O => \N__51393\,
            I => \N__51374\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__51390\,
            I => \N__51371\
        );

    \I__12303\ : Span4Mux_v
    port map (
            O => \N__51387\,
            I => \N__51368\
        );

    \I__12302\ : InMux
    port map (
            O => \N__51384\,
            I => \N__51365\
        );

    \I__12301\ : InMux
    port map (
            O => \N__51383\,
            I => \N__51362\
        );

    \I__12300\ : Span4Mux_v
    port map (
            O => \N__51380\,
            I => \N__51359\
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__51377\,
            I => \N__51356\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__51374\,
            I => \N__51353\
        );

    \I__12297\ : Span4Mux_v
    port map (
            O => \N__51371\,
            I => \N__51350\
        );

    \I__12296\ : Span4Mux_h
    port map (
            O => \N__51368\,
            I => \N__51343\
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__51365\,
            I => \N__51343\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__51362\,
            I => \N__51343\
        );

    \I__12293\ : Span4Mux_h
    port map (
            O => \N__51359\,
            I => \N__51335\
        );

    \I__12292\ : Span4Mux_v
    port map (
            O => \N__51356\,
            I => \N__51335\
        );

    \I__12291\ : Span4Mux_h
    port map (
            O => \N__51353\,
            I => \N__51335\
        );

    \I__12290\ : Span4Mux_v
    port map (
            O => \N__51350\,
            I => \N__51330\
        );

    \I__12289\ : Span4Mux_v
    port map (
            O => \N__51343\,
            I => \N__51330\
        );

    \I__12288\ : InMux
    port map (
            O => \N__51342\,
            I => \N__51327\
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__51335\,
            I => comm_rx_buf_7
        );

    \I__12286\ : Odrv4
    port map (
            O => \N__51330\,
            I => comm_rx_buf_7
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__51327\,
            I => comm_rx_buf_7
        );

    \I__12284\ : InMux
    port map (
            O => \N__51320\,
            I => \N__51314\
        );

    \I__12283\ : InMux
    port map (
            O => \N__51319\,
            I => \N__51314\
        );

    \I__12282\ : LocalMux
    port map (
            O => \N__51314\,
            I => \N__51308\
        );

    \I__12281\ : InMux
    port map (
            O => \N__51313\,
            I => \N__51303\
        );

    \I__12280\ : InMux
    port map (
            O => \N__51312\,
            I => \N__51303\
        );

    \I__12279\ : InMux
    port map (
            O => \N__51311\,
            I => \N__51300\
        );

    \I__12278\ : Span4Mux_h
    port map (
            O => \N__51308\,
            I => \N__51293\
        );

    \I__12277\ : LocalMux
    port map (
            O => \N__51303\,
            I => \N__51293\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__51300\,
            I => \N__51290\
        );

    \I__12275\ : InMux
    port map (
            O => \N__51299\,
            I => \N__51285\
        );

    \I__12274\ : InMux
    port map (
            O => \N__51298\,
            I => \N__51285\
        );

    \I__12273\ : Span4Mux_h
    port map (
            O => \N__51293\,
            I => \N__51281\
        );

    \I__12272\ : Span4Mux_v
    port map (
            O => \N__51290\,
            I => \N__51276\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__51285\,
            I => \N__51276\
        );

    \I__12270\ : InMux
    port map (
            O => \N__51284\,
            I => \N__51273\
        );

    \I__12269\ : Odrv4
    port map (
            O => \N__51281\,
            I => n12244
        );

    \I__12268\ : Odrv4
    port map (
            O => \N__51276\,
            I => n12244
        );

    \I__12267\ : LocalMux
    port map (
            O => \N__51273\,
            I => n12244
        );

    \I__12266\ : InMux
    port map (
            O => \N__51266\,
            I => \N__51262\
        );

    \I__12265\ : InMux
    port map (
            O => \N__51265\,
            I => \N__51259\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__51262\,
            I => comm_buf_6_7
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__51259\,
            I => comm_buf_6_7
        );

    \I__12262\ : InMux
    port map (
            O => \N__51254\,
            I => \N__51251\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__51251\,
            I => \N__51248\
        );

    \I__12260\ : Span4Mux_v
    port map (
            O => \N__51248\,
            I => \N__51245\
        );

    \I__12259\ : Span4Mux_v
    port map (
            O => \N__51245\,
            I => \N__51242\
        );

    \I__12258\ : Sp12to4
    port map (
            O => \N__51242\,
            I => \N__51239\
        );

    \I__12257\ : Span12Mux_h
    port map (
            O => \N__51239\,
            I => \N__51236\
        );

    \I__12256\ : Odrv12
    port map (
            O => \N__51236\,
            I => \THERMOSTAT\
        );

    \I__12255\ : InMux
    port map (
            O => \N__51233\,
            I => \N__51230\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__51230\,
            I => \N__51227\
        );

    \I__12253\ : Odrv4
    port map (
            O => \N__51227\,
            I => buf_control_7
        );

    \I__12252\ : CEMux
    port map (
            O => \N__51224\,
            I => \N__51221\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__51221\,
            I => \N__51218\
        );

    \I__12250\ : Span4Mux_v
    port map (
            O => \N__51218\,
            I => \N__51215\
        );

    \I__12249\ : Odrv4
    port map (
            O => \N__51215\,
            I => n11935
        );

    \I__12248\ : SRMux
    port map (
            O => \N__51212\,
            I => \N__51209\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__51209\,
            I => \N__51205\
        );

    \I__12246\ : SRMux
    port map (
            O => \N__51208\,
            I => \N__51202\
        );

    \I__12245\ : Span4Mux_v
    port map (
            O => \N__51205\,
            I => \N__51197\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__51202\,
            I => \N__51197\
        );

    \I__12243\ : Span4Mux_h
    port map (
            O => \N__51197\,
            I => \N__51194\
        );

    \I__12242\ : Span4Mux_h
    port map (
            O => \N__51194\,
            I => \N__51191\
        );

    \I__12241\ : Odrv4
    port map (
            O => \N__51191\,
            I => n19904
        );

    \I__12240\ : CascadeMux
    port map (
            O => \N__51188\,
            I => \N__51184\
        );

    \I__12239\ : CascadeMux
    port map (
            O => \N__51187\,
            I => \N__51178\
        );

    \I__12238\ : InMux
    port map (
            O => \N__51184\,
            I => \N__51175\
        );

    \I__12237\ : InMux
    port map (
            O => \N__51183\,
            I => \N__51172\
        );

    \I__12236\ : InMux
    port map (
            O => \N__51182\,
            I => \N__51169\
        );

    \I__12235\ : InMux
    port map (
            O => \N__51181\,
            I => \N__51165\
        );

    \I__12234\ : InMux
    port map (
            O => \N__51178\,
            I => \N__51162\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__51175\,
            I => \N__51157\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__51172\,
            I => \N__51157\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__51169\,
            I => \N__51154\
        );

    \I__12230\ : InMux
    port map (
            O => \N__51168\,
            I => \N__51151\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__51165\,
            I => \N__51148\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__51162\,
            I => \N__51145\
        );

    \I__12227\ : Span4Mux_v
    port map (
            O => \N__51157\,
            I => \N__51142\
        );

    \I__12226\ : Span4Mux_v
    port map (
            O => \N__51154\,
            I => \N__51139\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__51151\,
            I => \N__51136\
        );

    \I__12224\ : Span4Mux_v
    port map (
            O => \N__51148\,
            I => \N__51133\
        );

    \I__12223\ : Span4Mux_v
    port map (
            O => \N__51145\,
            I => \N__51124\
        );

    \I__12222\ : Span4Mux_h
    port map (
            O => \N__51142\,
            I => \N__51124\
        );

    \I__12221\ : Span4Mux_v
    port map (
            O => \N__51139\,
            I => \N__51124\
        );

    \I__12220\ : Span4Mux_v
    port map (
            O => \N__51136\,
            I => \N__51124\
        );

    \I__12219\ : Odrv4
    port map (
            O => \N__51133\,
            I => comm_buf_1_4
        );

    \I__12218\ : Odrv4
    port map (
            O => \N__51124\,
            I => comm_buf_1_4
        );

    \I__12217\ : InMux
    port map (
            O => \N__51119\,
            I => \N__51115\
        );

    \I__12216\ : InMux
    port map (
            O => \N__51118\,
            I => \N__51112\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__51115\,
            I => \N__51109\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__51112\,
            I => \N__51106\
        );

    \I__12213\ : Span4Mux_h
    port map (
            O => \N__51109\,
            I => \N__51103\
        );

    \I__12212\ : Span4Mux_h
    port map (
            O => \N__51106\,
            I => \N__51100\
        );

    \I__12211\ : Odrv4
    port map (
            O => \N__51103\,
            I => n14_adj_1548
        );

    \I__12210\ : Odrv4
    port map (
            O => \N__51100\,
            I => n14_adj_1548
        );

    \I__12209\ : InMux
    port map (
            O => \N__51095\,
            I => \N__51091\
        );

    \I__12208\ : CascadeMux
    port map (
            O => \N__51094\,
            I => \N__51088\
        );

    \I__12207\ : LocalMux
    port map (
            O => \N__51091\,
            I => \N__51085\
        );

    \I__12206\ : InMux
    port map (
            O => \N__51088\,
            I => \N__51082\
        );

    \I__12205\ : Span4Mux_v
    port map (
            O => \N__51085\,
            I => \N__51077\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__51082\,
            I => \N__51077\
        );

    \I__12203\ : Span4Mux_h
    port map (
            O => \N__51077\,
            I => \N__51073\
        );

    \I__12202\ : CascadeMux
    port map (
            O => \N__51076\,
            I => \N__51070\
        );

    \I__12201\ : Span4Mux_h
    port map (
            O => \N__51073\,
            I => \N__51067\
        );

    \I__12200\ : InMux
    port map (
            O => \N__51070\,
            I => \N__51064\
        );

    \I__12199\ : Odrv4
    port map (
            O => \N__51067\,
            I => cmd_rdadctmp_20_adj_1430
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__51064\,
            I => cmd_rdadctmp_20_adj_1430
        );

    \I__12197\ : CascadeMux
    port map (
            O => \N__51059\,
            I => \N__51056\
        );

    \I__12196\ : InMux
    port map (
            O => \N__51056\,
            I => \N__51051\
        );

    \I__12195\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51048\
        );

    \I__12194\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51044\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__51051\,
            I => \N__51039\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__51048\,
            I => \N__51036\
        );

    \I__12191\ : CascadeMux
    port map (
            O => \N__51047\,
            I => \N__51033\
        );

    \I__12190\ : LocalMux
    port map (
            O => \N__51044\,
            I => \N__51029\
        );

    \I__12189\ : InMux
    port map (
            O => \N__51043\,
            I => \N__51026\
        );

    \I__12188\ : InMux
    port map (
            O => \N__51042\,
            I => \N__51023\
        );

    \I__12187\ : Span4Mux_v
    port map (
            O => \N__51039\,
            I => \N__51018\
        );

    \I__12186\ : Span4Mux_v
    port map (
            O => \N__51036\,
            I => \N__51018\
        );

    \I__12185\ : InMux
    port map (
            O => \N__51033\,
            I => \N__51015\
        );

    \I__12184\ : InMux
    port map (
            O => \N__51032\,
            I => \N__51012\
        );

    \I__12183\ : Span4Mux_v
    port map (
            O => \N__51029\,
            I => \N__51009\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__51026\,
            I => \N__51006\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__51023\,
            I => \N__51003\
        );

    \I__12180\ : Span4Mux_h
    port map (
            O => \N__51018\,
            I => \N__50996\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__51015\,
            I => \N__50996\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__51012\,
            I => \N__50996\
        );

    \I__12177\ : Span4Mux_v
    port map (
            O => \N__51009\,
            I => \N__50989\
        );

    \I__12176\ : Span4Mux_h
    port map (
            O => \N__51006\,
            I => \N__50989\
        );

    \I__12175\ : Span4Mux_v
    port map (
            O => \N__51003\,
            I => \N__50984\
        );

    \I__12174\ : Span4Mux_v
    port map (
            O => \N__50996\,
            I => \N__50984\
        );

    \I__12173\ : InMux
    port map (
            O => \N__50995\,
            I => \N__50981\
        );

    \I__12172\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50978\
        );

    \I__12171\ : Odrv4
    port map (
            O => \N__50989\,
            I => comm_rx_buf_5
        );

    \I__12170\ : Odrv4
    port map (
            O => \N__50984\,
            I => comm_rx_buf_5
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__50981\,
            I => comm_rx_buf_5
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__50978\,
            I => comm_rx_buf_5
        );

    \I__12167\ : CascadeMux
    port map (
            O => \N__50969\,
            I => \N__50965\
        );

    \I__12166\ : InMux
    port map (
            O => \N__50968\,
            I => \N__50960\
        );

    \I__12165\ : InMux
    port map (
            O => \N__50965\,
            I => \N__50960\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__50960\,
            I => comm_buf_6_5
        );

    \I__12163\ : CascadeMux
    port map (
            O => \N__50957\,
            I => \n2369_cascade_\
        );

    \I__12162\ : CascadeMux
    port map (
            O => \N__50954\,
            I => \n21130_cascade_\
        );

    \I__12161\ : CEMux
    port map (
            O => \N__50951\,
            I => \N__50948\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__50948\,
            I => \N__50945\
        );

    \I__12159\ : Odrv4
    port map (
            O => \N__50945\,
            I => n14_adj_1506
        );

    \I__12158\ : InMux
    port map (
            O => \N__50942\,
            I => \N__50939\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__50939\,
            I => \N__50936\
        );

    \I__12156\ : Odrv4
    port map (
            O => \N__50936\,
            I => n3
        );

    \I__12155\ : CascadeMux
    port map (
            O => \N__50933\,
            I => \N__50927\
        );

    \I__12154\ : InMux
    port map (
            O => \N__50932\,
            I => \N__50922\
        );

    \I__12153\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50917\
        );

    \I__12152\ : InMux
    port map (
            O => \N__50930\,
            I => \N__50917\
        );

    \I__12151\ : InMux
    port map (
            O => \N__50927\,
            I => \N__50914\
        );

    \I__12150\ : InMux
    port map (
            O => \N__50926\,
            I => \N__50911\
        );

    \I__12149\ : InMux
    port map (
            O => \N__50925\,
            I => \N__50908\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__50922\,
            I => \N__50903\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__50917\,
            I => \N__50898\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__50914\,
            I => \N__50898\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__50911\,
            I => \N__50895\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__50908\,
            I => \N__50892\
        );

    \I__12143\ : InMux
    port map (
            O => \N__50907\,
            I => \N__50887\
        );

    \I__12142\ : InMux
    port map (
            O => \N__50906\,
            I => \N__50887\
        );

    \I__12141\ : Span4Mux_h
    port map (
            O => \N__50903\,
            I => \N__50882\
        );

    \I__12140\ : Span4Mux_v
    port map (
            O => \N__50898\,
            I => \N__50879\
        );

    \I__12139\ : Span4Mux_h
    port map (
            O => \N__50895\,
            I => \N__50872\
        );

    \I__12138\ : Span4Mux_h
    port map (
            O => \N__50892\,
            I => \N__50872\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__50887\,
            I => \N__50872\
        );

    \I__12136\ : InMux
    port map (
            O => \N__50886\,
            I => \N__50867\
        );

    \I__12135\ : InMux
    port map (
            O => \N__50885\,
            I => \N__50867\
        );

    \I__12134\ : Odrv4
    port map (
            O => \N__50882\,
            I => n20681
        );

    \I__12133\ : Odrv4
    port map (
            O => \N__50879\,
            I => n20681
        );

    \I__12132\ : Odrv4
    port map (
            O => \N__50872\,
            I => n20681
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__50867\,
            I => n20681
        );

    \I__12130\ : CascadeMux
    port map (
            O => \N__50858\,
            I => \n3_cascade_\
        );

    \I__12129\ : InMux
    port map (
            O => \N__50855\,
            I => \N__50851\
        );

    \I__12128\ : InMux
    port map (
            O => \N__50854\,
            I => \N__50847\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__50851\,
            I => \N__50844\
        );

    \I__12126\ : InMux
    port map (
            O => \N__50850\,
            I => \N__50841\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__50847\,
            I => n2369
        );

    \I__12124\ : Odrv4
    port map (
            O => \N__50844\,
            I => n2369
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__50841\,
            I => n2369
        );

    \I__12122\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50831\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__50831\,
            I => n19655
        );

    \I__12120\ : InMux
    port map (
            O => \N__50828\,
            I => \N__50825\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__50825\,
            I => n23_adj_1501
        );

    \I__12118\ : CascadeMux
    port map (
            O => \N__50822\,
            I => \n21_adj_1600_cascade_\
        );

    \I__12117\ : InMux
    port map (
            O => \N__50819\,
            I => \N__50816\
        );

    \I__12116\ : LocalMux
    port map (
            O => \N__50816\,
            I => n17485
        );

    \I__12115\ : CEMux
    port map (
            O => \N__50813\,
            I => \N__50810\
        );

    \I__12114\ : LocalMux
    port map (
            O => \N__50810\,
            I => \N__50807\
        );

    \I__12113\ : Odrv12
    port map (
            O => \N__50807\,
            I => n18_adj_1633
        );

    \I__12112\ : CascadeMux
    port map (
            O => \N__50804\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50801\,
            I => \N__50798\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__50798\,
            I => \comm_spi.n22667\
        );

    \I__12109\ : InMux
    port map (
            O => \N__50795\,
            I => \N__50792\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__50792\,
            I => \N__50789\
        );

    \I__12107\ : Odrv4
    port map (
            O => \N__50789\,
            I => \comm_spi.n14630\
        );

    \I__12106\ : CascadeMux
    port map (
            O => \N__50786\,
            I => \comm_spi.n22667_cascade_\
        );

    \I__12105\ : InMux
    port map (
            O => \N__50783\,
            I => \N__50779\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50782\,
            I => \N__50772\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__50779\,
            I => \N__50768\
        );

    \I__12102\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50765\
        );

    \I__12101\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50762\
        );

    \I__12100\ : InMux
    port map (
            O => \N__50776\,
            I => \N__50758\
        );

    \I__12099\ : InMux
    port map (
            O => \N__50775\,
            I => \N__50755\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__50772\,
            I => \N__50752\
        );

    \I__12097\ : InMux
    port map (
            O => \N__50771\,
            I => \N__50749\
        );

    \I__12096\ : Span4Mux_h
    port map (
            O => \N__50768\,
            I => \N__50742\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__50765\,
            I => \N__50742\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__50762\,
            I => \N__50742\
        );

    \I__12093\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50739\
        );

    \I__12092\ : LocalMux
    port map (
            O => \N__50758\,
            I => \N__50736\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__50755\,
            I => \N__50733\
        );

    \I__12090\ : Span4Mux_v
    port map (
            O => \N__50752\,
            I => \N__50728\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__50749\,
            I => \N__50728\
        );

    \I__12088\ : Span4Mux_v
    port map (
            O => \N__50742\,
            I => \N__50723\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__50739\,
            I => \N__50723\
        );

    \I__12086\ : Span12Mux_h
    port map (
            O => \N__50736\,
            I => \N__50720\
        );

    \I__12085\ : Span4Mux_v
    port map (
            O => \N__50733\,
            I => \N__50715\
        );

    \I__12084\ : Span4Mux_v
    port map (
            O => \N__50728\,
            I => \N__50715\
        );

    \I__12083\ : Span4Mux_h
    port map (
            O => \N__50723\,
            I => \N__50712\
        );

    \I__12082\ : Odrv12
    port map (
            O => \N__50720\,
            I => comm_rx_buf_0
        );

    \I__12081\ : Odrv4
    port map (
            O => \N__50715\,
            I => comm_rx_buf_0
        );

    \I__12080\ : Odrv4
    port map (
            O => \N__50712\,
            I => comm_rx_buf_0
        );

    \I__12079\ : CascadeMux
    port map (
            O => \N__50705\,
            I => \comm_rx_buf_0_cascade_\
        );

    \I__12078\ : InMux
    port map (
            O => \N__50702\,
            I => \N__50698\
        );

    \I__12077\ : InMux
    port map (
            O => \N__50701\,
            I => \N__50695\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__50698\,
            I => \N__50692\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__50695\,
            I => comm_buf_6_0
        );

    \I__12074\ : Odrv12
    port map (
            O => \N__50692\,
            I => comm_buf_6_0
        );

    \I__12073\ : InMux
    port map (
            O => \N__50687\,
            I => \N__50671\
        );

    \I__12072\ : InMux
    port map (
            O => \N__50686\,
            I => \N__50671\
        );

    \I__12071\ : InMux
    port map (
            O => \N__50685\,
            I => \N__50671\
        );

    \I__12070\ : InMux
    port map (
            O => \N__50684\,
            I => \N__50659\
        );

    \I__12069\ : InMux
    port map (
            O => \N__50683\,
            I => \N__50652\
        );

    \I__12068\ : InMux
    port map (
            O => \N__50682\,
            I => \N__50652\
        );

    \I__12067\ : InMux
    port map (
            O => \N__50681\,
            I => \N__50652\
        );

    \I__12066\ : InMux
    port map (
            O => \N__50680\,
            I => \N__50645\
        );

    \I__12065\ : InMux
    port map (
            O => \N__50679\,
            I => \N__50645\
        );

    \I__12064\ : InMux
    port map (
            O => \N__50678\,
            I => \N__50645\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__50671\,
            I => \N__50642\
        );

    \I__12062\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50637\
        );

    \I__12061\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50637\
        );

    \I__12060\ : CascadeMux
    port map (
            O => \N__50668\,
            I => \N__50633\
        );

    \I__12059\ : InMux
    port map (
            O => \N__50667\,
            I => \N__50626\
        );

    \I__12058\ : InMux
    port map (
            O => \N__50666\,
            I => \N__50626\
        );

    \I__12057\ : InMux
    port map (
            O => \N__50665\,
            I => \N__50619\
        );

    \I__12056\ : InMux
    port map (
            O => \N__50664\,
            I => \N__50619\
        );

    \I__12055\ : InMux
    port map (
            O => \N__50663\,
            I => \N__50619\
        );

    \I__12054\ : InMux
    port map (
            O => \N__50662\,
            I => \N__50616\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__50659\,
            I => \N__50613\
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__50652\,
            I => \N__50604\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__50645\,
            I => \N__50604\
        );

    \I__12050\ : Span4Mux_v
    port map (
            O => \N__50642\,
            I => \N__50604\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__50637\,
            I => \N__50604\
        );

    \I__12048\ : InMux
    port map (
            O => \N__50636\,
            I => \N__50601\
        );

    \I__12047\ : InMux
    port map (
            O => \N__50633\,
            I => \N__50598\
        );

    \I__12046\ : InMux
    port map (
            O => \N__50632\,
            I => \N__50593\
        );

    \I__12045\ : InMux
    port map (
            O => \N__50631\,
            I => \N__50593\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__50626\,
            I => \N__50590\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__50619\,
            I => \N__50585\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__50616\,
            I => \N__50585\
        );

    \I__12041\ : Span4Mux_v
    port map (
            O => \N__50613\,
            I => \N__50580\
        );

    \I__12040\ : Span4Mux_h
    port map (
            O => \N__50604\,
            I => \N__50580\
        );

    \I__12039\ : LocalMux
    port map (
            O => \N__50601\,
            I => comm_index_2
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__50598\,
            I => comm_index_2
        );

    \I__12037\ : LocalMux
    port map (
            O => \N__50593\,
            I => comm_index_2
        );

    \I__12036\ : Odrv4
    port map (
            O => \N__50590\,
            I => comm_index_2
        );

    \I__12035\ : Odrv4
    port map (
            O => \N__50585\,
            I => comm_index_2
        );

    \I__12034\ : Odrv4
    port map (
            O => \N__50580\,
            I => comm_index_2
        );

    \I__12033\ : InMux
    port map (
            O => \N__50567\,
            I => \N__50564\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__50564\,
            I => \N__50561\
        );

    \I__12031\ : Span4Mux_h
    port map (
            O => \N__50561\,
            I => \N__50558\
        );

    \I__12030\ : Odrv4
    port map (
            O => \N__50558\,
            I => comm_buf_2_5
        );

    \I__12029\ : CascadeMux
    port map (
            O => \N__50555\,
            I => \N__50549\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50539\
        );

    \I__12027\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50539\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50529\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50549\,
            I => \N__50526\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50548\,
            I => \N__50523\
        );

    \I__12023\ : InMux
    port map (
            O => \N__50547\,
            I => \N__50518\
        );

    \I__12022\ : InMux
    port map (
            O => \N__50546\,
            I => \N__50518\
        );

    \I__12021\ : InMux
    port map (
            O => \N__50545\,
            I => \N__50513\
        );

    \I__12020\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50513\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__50539\,
            I => \N__50510\
        );

    \I__12018\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50507\
        );

    \I__12017\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50499\
        );

    \I__12016\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50499\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50535\,
            I => \N__50499\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50534\,
            I => \N__50496\
        );

    \I__12013\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50488\
        );

    \I__12012\ : InMux
    port map (
            O => \N__50532\,
            I => \N__50488\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__50529\,
            I => \N__50485\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__50526\,
            I => \N__50478\
        );

    \I__12009\ : LocalMux
    port map (
            O => \N__50523\,
            I => \N__50475\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__50518\,
            I => \N__50466\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__50513\,
            I => \N__50466\
        );

    \I__12006\ : Span4Mux_v
    port map (
            O => \N__50510\,
            I => \N__50466\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__50507\,
            I => \N__50466\
        );

    \I__12004\ : InMux
    port map (
            O => \N__50506\,
            I => \N__50463\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50458\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50496\,
            I => \N__50458\
        );

    \I__12001\ : InMux
    port map (
            O => \N__50495\,
            I => \N__50451\
        );

    \I__12000\ : InMux
    port map (
            O => \N__50494\,
            I => \N__50451\
        );

    \I__11999\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50451\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50488\,
            I => \N__50448\
        );

    \I__11997\ : Span4Mux_h
    port map (
            O => \N__50485\,
            I => \N__50445\
        );

    \I__11996\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50436\
        );

    \I__11995\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50436\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50482\,
            I => \N__50436\
        );

    \I__11993\ : InMux
    port map (
            O => \N__50481\,
            I => \N__50436\
        );

    \I__11992\ : Span4Mux_h
    port map (
            O => \N__50478\,
            I => \N__50429\
        );

    \I__11991\ : Span4Mux_h
    port map (
            O => \N__50475\,
            I => \N__50429\
        );

    \I__11990\ : Span4Mux_h
    port map (
            O => \N__50466\,
            I => \N__50429\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__50463\,
            I => comm_index_1
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__50458\,
            I => comm_index_1
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__50451\,
            I => comm_index_1
        );

    \I__11986\ : Odrv12
    port map (
            O => \N__50448\,
            I => comm_index_1
        );

    \I__11985\ : Odrv4
    port map (
            O => \N__50445\,
            I => comm_index_1
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__50436\,
            I => comm_index_1
        );

    \I__11983\ : Odrv4
    port map (
            O => \N__50429\,
            I => comm_index_1
        );

    \I__11982\ : InMux
    port map (
            O => \N__50414\,
            I => \N__50411\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__50411\,
            I => \N__50408\
        );

    \I__11980\ : Odrv12
    port map (
            O => \N__50408\,
            I => n22172
        );

    \I__11979\ : SRMux
    port map (
            O => \N__50405\,
            I => \N__50402\
        );

    \I__11978\ : LocalMux
    port map (
            O => \N__50402\,
            I => \N__50399\
        );

    \I__11977\ : Odrv4
    port map (
            O => \N__50399\,
            I => n14671
        );

    \I__11976\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50393\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__50393\,
            I => \SIG_DDS.n21331\
        );

    \I__11974\ : CascadeMux
    port map (
            O => \N__50390\,
            I => \N__50387\
        );

    \I__11973\ : InMux
    port map (
            O => \N__50387\,
            I => \N__50384\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__50384\,
            I => \SIG_DDS.n10\
        );

    \I__11971\ : CEMux
    port map (
            O => \N__50381\,
            I => \N__50377\
        );

    \I__11970\ : CEMux
    port map (
            O => \N__50380\,
            I => \N__50374\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__50377\,
            I => \N__50371\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__50374\,
            I => \SIG_DDS.n9\
        );

    \I__11967\ : Odrv4
    port map (
            O => \N__50371\,
            I => \SIG_DDS.n9\
        );

    \I__11966\ : InMux
    port map (
            O => \N__50366\,
            I => \N__50363\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__50363\,
            I => \N__50355\
        );

    \I__11964\ : CascadeMux
    port map (
            O => \N__50362\,
            I => \N__50350\
        );

    \I__11963\ : InMux
    port map (
            O => \N__50361\,
            I => \N__50346\
        );

    \I__11962\ : InMux
    port map (
            O => \N__50360\,
            I => \N__50343\
        );

    \I__11961\ : InMux
    port map (
            O => \N__50359\,
            I => \N__50340\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50358\,
            I => \N__50337\
        );

    \I__11959\ : Span12Mux_s8_v
    port map (
            O => \N__50355\,
            I => \N__50334\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50329\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50353\,
            I => \N__50329\
        );

    \I__11956\ : InMux
    port map (
            O => \N__50350\,
            I => \N__50324\
        );

    \I__11955\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50324\
        );

    \I__11954\ : LocalMux
    port map (
            O => \N__50346\,
            I => dds_state_0
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__50343\,
            I => dds_state_0
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__50340\,
            I => dds_state_0
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__50337\,
            I => dds_state_0
        );

    \I__11950\ : Odrv12
    port map (
            O => \N__50334\,
            I => dds_state_0
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__50329\,
            I => dds_state_0
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__50324\,
            I => dds_state_0
        );

    \I__11947\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50278\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50308\,
            I => \N__50278\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50278\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50278\
        );

    \I__11943\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50278\
        );

    \I__11942\ : InMux
    port map (
            O => \N__50304\,
            I => \N__50278\
        );

    \I__11941\ : InMux
    port map (
            O => \N__50303\,
            I => \N__50278\
        );

    \I__11940\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50278\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50263\
        );

    \I__11938\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50263\
        );

    \I__11937\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50263\
        );

    \I__11936\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50263\
        );

    \I__11935\ : InMux
    port map (
            O => \N__50297\,
            I => \N__50263\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50296\,
            I => \N__50263\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50295\,
            I => \N__50263\
        );

    \I__11932\ : LocalMux
    port map (
            O => \N__50278\,
            I => \N__50255\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__50263\,
            I => \N__50255\
        );

    \I__11930\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50251\
        );

    \I__11929\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50243\
        );

    \I__11928\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50243\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__50255\,
            I => \N__50240\
        );

    \I__11926\ : InMux
    port map (
            O => \N__50254\,
            I => \N__50237\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__50251\,
            I => \N__50234\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50250\,
            I => \N__50230\
        );

    \I__11923\ : InMux
    port map (
            O => \N__50249\,
            I => \N__50225\
        );

    \I__11922\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50225\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__50243\,
            I => \N__50220\
        );

    \I__11920\ : Span4Mux_h
    port map (
            O => \N__50240\,
            I => \N__50213\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__50237\,
            I => \N__50213\
        );

    \I__11918\ : Span4Mux_v
    port map (
            O => \N__50234\,
            I => \N__50213\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50210\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__50230\,
            I => \N__50205\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__50225\,
            I => \N__50205\
        );

    \I__11914\ : InMux
    port map (
            O => \N__50224\,
            I => \N__50200\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50223\,
            I => \N__50200\
        );

    \I__11912\ : Span4Mux_v
    port map (
            O => \N__50220\,
            I => \N__50197\
        );

    \I__11911\ : Odrv4
    port map (
            O => \N__50213\,
            I => dds_state_2
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__50210\,
            I => dds_state_2
        );

    \I__11909\ : Odrv12
    port map (
            O => \N__50205\,
            I => dds_state_2
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__50200\,
            I => dds_state_2
        );

    \I__11907\ : Odrv4
    port map (
            O => \N__50197\,
            I => dds_state_2
        );

    \I__11906\ : SRMux
    port map (
            O => \N__50186\,
            I => \N__50173\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50185\,
            I => \N__50158\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50184\,
            I => \N__50158\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50183\,
            I => \N__50158\
        );

    \I__11902\ : InMux
    port map (
            O => \N__50182\,
            I => \N__50158\
        );

    \I__11901\ : InMux
    port map (
            O => \N__50181\,
            I => \N__50158\
        );

    \I__11900\ : InMux
    port map (
            O => \N__50180\,
            I => \N__50158\
        );

    \I__11899\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50158\
        );

    \I__11898\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50151\
        );

    \I__11897\ : InMux
    port map (
            O => \N__50177\,
            I => \N__50151\
        );

    \I__11896\ : CEMux
    port map (
            O => \N__50176\,
            I => \N__50148\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__50173\,
            I => \N__50145\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50158\,
            I => \N__50142\
        );

    \I__11893\ : CascadeMux
    port map (
            O => \N__50157\,
            I => \N__50134\
        );

    \I__11892\ : InMux
    port map (
            O => \N__50156\,
            I => \N__50127\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__50151\,
            I => \N__50124\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__50148\,
            I => \N__50121\
        );

    \I__11889\ : Span4Mux_v
    port map (
            O => \N__50145\,
            I => \N__50116\
        );

    \I__11888\ : Span4Mux_h
    port map (
            O => \N__50142\,
            I => \N__50116\
        );

    \I__11887\ : InMux
    port map (
            O => \N__50141\,
            I => \N__50099\
        );

    \I__11886\ : InMux
    port map (
            O => \N__50140\,
            I => \N__50099\
        );

    \I__11885\ : InMux
    port map (
            O => \N__50139\,
            I => \N__50099\
        );

    \I__11884\ : InMux
    port map (
            O => \N__50138\,
            I => \N__50099\
        );

    \I__11883\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50099\
        );

    \I__11882\ : InMux
    port map (
            O => \N__50134\,
            I => \N__50099\
        );

    \I__11881\ : InMux
    port map (
            O => \N__50133\,
            I => \N__50099\
        );

    \I__11880\ : InMux
    port map (
            O => \N__50132\,
            I => \N__50099\
        );

    \I__11879\ : InMux
    port map (
            O => \N__50131\,
            I => \N__50095\
        );

    \I__11878\ : InMux
    port map (
            O => \N__50130\,
            I => \N__50092\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__50127\,
            I => \N__50087\
        );

    \I__11876\ : Span4Mux_h
    port map (
            O => \N__50124\,
            I => \N__50087\
        );

    \I__11875\ : Span4Mux_h
    port map (
            O => \N__50121\,
            I => \N__50077\
        );

    \I__11874\ : Span4Mux_h
    port map (
            O => \N__50116\,
            I => \N__50077\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__50099\,
            I => \N__50074\
        );

    \I__11872\ : InMux
    port map (
            O => \N__50098\,
            I => \N__50071\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__50095\,
            I => \N__50064\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__50092\,
            I => \N__50064\
        );

    \I__11869\ : Span4Mux_h
    port map (
            O => \N__50087\,
            I => \N__50064\
        );

    \I__11868\ : InMux
    port map (
            O => \N__50086\,
            I => \N__50057\
        );

    \I__11867\ : InMux
    port map (
            O => \N__50085\,
            I => \N__50057\
        );

    \I__11866\ : InMux
    port map (
            O => \N__50084\,
            I => \N__50057\
        );

    \I__11865\ : InMux
    port map (
            O => \N__50083\,
            I => \N__50052\
        );

    \I__11864\ : InMux
    port map (
            O => \N__50082\,
            I => \N__50052\
        );

    \I__11863\ : Odrv4
    port map (
            O => \N__50077\,
            I => dds_state_1
        );

    \I__11862\ : Odrv12
    port map (
            O => \N__50074\,
            I => dds_state_1
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__50071\,
            I => dds_state_1
        );

    \I__11860\ : Odrv4
    port map (
            O => \N__50064\,
            I => dds_state_1
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__50057\,
            I => dds_state_1
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__50052\,
            I => dds_state_1
        );

    \I__11857\ : IoInMux
    port map (
            O => \N__50039\,
            I => \N__50036\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__50036\,
            I => \N__50033\
        );

    \I__11855\ : IoSpan4Mux
    port map (
            O => \N__50033\,
            I => \N__50030\
        );

    \I__11854\ : IoSpan4Mux
    port map (
            O => \N__50030\,
            I => \N__50027\
        );

    \I__11853\ : Span4Mux_s3_v
    port map (
            O => \N__50027\,
            I => \N__50023\
        );

    \I__11852\ : CascadeMux
    port map (
            O => \N__50026\,
            I => \N__50020\
        );

    \I__11851\ : Span4Mux_v
    port map (
            O => \N__50023\,
            I => \N__50017\
        );

    \I__11850\ : InMux
    port map (
            O => \N__50020\,
            I => \N__50014\
        );

    \I__11849\ : Odrv4
    port map (
            O => \N__50017\,
            I => \DDS_SCK\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__50014\,
            I => \DDS_SCK\
        );

    \I__11847\ : InMux
    port map (
            O => \N__50009\,
            I => \N__50006\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__50006\,
            I => \N__50003\
        );

    \I__11845\ : Span4Mux_v
    port map (
            O => \N__50003\,
            I => \N__49999\
        );

    \I__11844\ : InMux
    port map (
            O => \N__50002\,
            I => \N__49995\
        );

    \I__11843\ : Sp12to4
    port map (
            O => \N__49999\,
            I => \N__49992\
        );

    \I__11842\ : InMux
    port map (
            O => \N__49998\,
            I => \N__49989\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__49995\,
            I => \N__49986\
        );

    \I__11840\ : Odrv12
    port map (
            O => \N__49992\,
            I => wdtick_flag
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__49989\,
            I => wdtick_flag
        );

    \I__11838\ : Odrv4
    port map (
            O => \N__49986\,
            I => wdtick_flag
        );

    \I__11837\ : InMux
    port map (
            O => \N__49979\,
            I => \N__49975\
        );

    \I__11836\ : InMux
    port map (
            O => \N__49978\,
            I => \N__49972\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__49975\,
            I => \N__49968\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__49972\,
            I => \N__49965\
        );

    \I__11833\ : InMux
    port map (
            O => \N__49971\,
            I => \N__49962\
        );

    \I__11832\ : Span4Mux_v
    port map (
            O => \N__49968\,
            I => \N__49959\
        );

    \I__11831\ : Odrv4
    port map (
            O => \N__49965\,
            I => buf_control_0
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__49962\,
            I => buf_control_0
        );

    \I__11829\ : Odrv4
    port map (
            O => \N__49959\,
            I => buf_control_0
        );

    \I__11828\ : IoInMux
    port map (
            O => \N__49952\,
            I => \N__49949\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49949\,
            I => \N__49946\
        );

    \I__11826\ : IoSpan4Mux
    port map (
            O => \N__49946\,
            I => \N__49943\
        );

    \I__11825\ : Span4Mux_s3_v
    port map (
            O => \N__49943\,
            I => \N__49940\
        );

    \I__11824\ : Span4Mux_v
    port map (
            O => \N__49940\,
            I => \N__49937\
        );

    \I__11823\ : Odrv4
    port map (
            O => \N__49937\,
            I => \CONT_SD\
        );

    \I__11822\ : InMux
    port map (
            O => \N__49934\,
            I => \N__49931\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__49931\,
            I => \N__49928\
        );

    \I__11820\ : Odrv4
    port map (
            O => \N__49928\,
            I => n20608
        );

    \I__11819\ : CascadeMux
    port map (
            O => \N__49925\,
            I => \N__49911\
        );

    \I__11818\ : CascadeMux
    port map (
            O => \N__49924\,
            I => \N__49905\
        );

    \I__11817\ : CascadeMux
    port map (
            O => \N__49923\,
            I => \N__49901\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49922\,
            I => \N__49890\
        );

    \I__11815\ : InMux
    port map (
            O => \N__49921\,
            I => \N__49890\
        );

    \I__11814\ : InMux
    port map (
            O => \N__49920\,
            I => \N__49887\
        );

    \I__11813\ : InMux
    port map (
            O => \N__49919\,
            I => \N__49882\
        );

    \I__11812\ : InMux
    port map (
            O => \N__49918\,
            I => \N__49882\
        );

    \I__11811\ : CascadeMux
    port map (
            O => \N__49917\,
            I => \N__49879\
        );

    \I__11810\ : CascadeMux
    port map (
            O => \N__49916\,
            I => \N__49876\
        );

    \I__11809\ : CascadeMux
    port map (
            O => \N__49915\,
            I => \N__49872\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49914\,
            I => \N__49868\
        );

    \I__11807\ : InMux
    port map (
            O => \N__49911\,
            I => \N__49861\
        );

    \I__11806\ : InMux
    port map (
            O => \N__49910\,
            I => \N__49861\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49909\,
            I => \N__49861\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49908\,
            I => \N__49856\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49905\,
            I => \N__49856\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49904\,
            I => \N__49849\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49901\,
            I => \N__49849\
        );

    \I__11800\ : InMux
    port map (
            O => \N__49900\,
            I => \N__49849\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49899\,
            I => \N__49840\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49898\,
            I => \N__49840\
        );

    \I__11797\ : InMux
    port map (
            O => \N__49897\,
            I => \N__49840\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49896\,
            I => \N__49840\
        );

    \I__11795\ : CascadeMux
    port map (
            O => \N__49895\,
            I => \N__49835\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49890\,
            I => \N__49820\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__49887\,
            I => \N__49815\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__49882\,
            I => \N__49815\
        );

    \I__11791\ : InMux
    port map (
            O => \N__49879\,
            I => \N__49810\
        );

    \I__11790\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49810\
        );

    \I__11789\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49803\
        );

    \I__11788\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49803\
        );

    \I__11787\ : InMux
    port map (
            O => \N__49871\,
            I => \N__49803\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__49868\,
            I => \N__49792\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__49861\,
            I => \N__49792\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__49856\,
            I => \N__49792\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__49849\,
            I => \N__49792\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49840\,
            I => \N__49792\
        );

    \I__11781\ : InMux
    port map (
            O => \N__49839\,
            I => \N__49785\
        );

    \I__11780\ : InMux
    port map (
            O => \N__49838\,
            I => \N__49785\
        );

    \I__11779\ : InMux
    port map (
            O => \N__49835\,
            I => \N__49785\
        );

    \I__11778\ : InMux
    port map (
            O => \N__49834\,
            I => \N__49782\
        );

    \I__11777\ : CascadeMux
    port map (
            O => \N__49833\,
            I => \N__49777\
        );

    \I__11776\ : CascadeMux
    port map (
            O => \N__49832\,
            I => \N__49768\
        );

    \I__11775\ : InMux
    port map (
            O => \N__49831\,
            I => \N__49762\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49762\
        );

    \I__11773\ : CascadeMux
    port map (
            O => \N__49829\,
            I => \N__49759\
        );

    \I__11772\ : InMux
    port map (
            O => \N__49828\,
            I => \N__49755\
        );

    \I__11771\ : CascadeMux
    port map (
            O => \N__49827\,
            I => \N__49751\
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__49826\,
            I => \N__49746\
        );

    \I__11769\ : CascadeMux
    port map (
            O => \N__49825\,
            I => \N__49743\
        );

    \I__11768\ : CascadeMux
    port map (
            O => \N__49824\,
            I => \N__49740\
        );

    \I__11767\ : CascadeMux
    port map (
            O => \N__49823\,
            I => \N__49736\
        );

    \I__11766\ : Span4Mux_h
    port map (
            O => \N__49820\,
            I => \N__49721\
        );

    \I__11765\ : Span4Mux_v
    port map (
            O => \N__49815\,
            I => \N__49721\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49810\,
            I => \N__49721\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__49803\,
            I => \N__49721\
        );

    \I__11762\ : Span4Mux_v
    port map (
            O => \N__49792\,
            I => \N__49721\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__49785\,
            I => \N__49721\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__49782\,
            I => \N__49717\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49714\
        );

    \I__11758\ : CascadeMux
    port map (
            O => \N__49780\,
            I => \N__49711\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49705\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49702\
        );

    \I__11755\ : CascadeMux
    port map (
            O => \N__49775\,
            I => \N__49695\
        );

    \I__11754\ : CascadeMux
    port map (
            O => \N__49774\,
            I => \N__49692\
        );

    \I__11753\ : CascadeMux
    port map (
            O => \N__49773\,
            I => \N__49688\
        );

    \I__11752\ : CascadeMux
    port map (
            O => \N__49772\,
            I => \N__49683\
        );

    \I__11751\ : CascadeMux
    port map (
            O => \N__49771\,
            I => \N__49679\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49674\
        );

    \I__11749\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49674\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49762\,
            I => \N__49671\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49759\,
            I => \N__49668\
        );

    \I__11746\ : CascadeMux
    port map (
            O => \N__49758\,
            I => \N__49665\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__49755\,
            I => \N__49660\
        );

    \I__11744\ : InMux
    port map (
            O => \N__49754\,
            I => \N__49657\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49652\
        );

    \I__11742\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49652\
        );

    \I__11741\ : InMux
    port map (
            O => \N__49749\,
            I => \N__49647\
        );

    \I__11740\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49647\
        );

    \I__11739\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49642\
        );

    \I__11738\ : InMux
    port map (
            O => \N__49740\,
            I => \N__49642\
        );

    \I__11737\ : InMux
    port map (
            O => \N__49739\,
            I => \N__49639\
        );

    \I__11736\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49631\
        );

    \I__11735\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49631\
        );

    \I__11734\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49631\
        );

    \I__11733\ : Span4Mux_v
    port map (
            O => \N__49721\,
            I => \N__49623\
        );

    \I__11732\ : InMux
    port map (
            O => \N__49720\,
            I => \N__49620\
        );

    \I__11731\ : Span4Mux_v
    port map (
            O => \N__49717\,
            I => \N__49617\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__49714\,
            I => \N__49614\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49711\,
            I => \N__49605\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49605\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49709\,
            I => \N__49605\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49708\,
            I => \N__49605\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__49705\,
            I => \N__49602\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__49702\,
            I => \N__49599\
        );

    \I__11723\ : CascadeMux
    port map (
            O => \N__49701\,
            I => \N__49596\
        );

    \I__11722\ : CascadeMux
    port map (
            O => \N__49700\,
            I => \N__49587\
        );

    \I__11721\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49576\
        );

    \I__11720\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49576\
        );

    \I__11719\ : InMux
    port map (
            O => \N__49695\,
            I => \N__49576\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49692\,
            I => \N__49576\
        );

    \I__11717\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49576\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49688\,
            I => \N__49569\
        );

    \I__11715\ : InMux
    port map (
            O => \N__49687\,
            I => \N__49569\
        );

    \I__11714\ : InMux
    port map (
            O => \N__49686\,
            I => \N__49569\
        );

    \I__11713\ : InMux
    port map (
            O => \N__49683\,
            I => \N__49562\
        );

    \I__11712\ : InMux
    port map (
            O => \N__49682\,
            I => \N__49562\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49679\,
            I => \N__49562\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__49674\,
            I => \N__49555\
        );

    \I__11709\ : Span4Mux_h
    port map (
            O => \N__49671\,
            I => \N__49555\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__49668\,
            I => \N__49555\
        );

    \I__11707\ : InMux
    port map (
            O => \N__49665\,
            I => \N__49548\
        );

    \I__11706\ : InMux
    port map (
            O => \N__49664\,
            I => \N__49548\
        );

    \I__11705\ : InMux
    port map (
            O => \N__49663\,
            I => \N__49548\
        );

    \I__11704\ : Span4Mux_v
    port map (
            O => \N__49660\,
            I => \N__49539\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__49657\,
            I => \N__49539\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__49652\,
            I => \N__49539\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__49647\,
            I => \N__49539\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__49642\,
            I => \N__49536\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__49639\,
            I => \N__49533\
        );

    \I__11698\ : InMux
    port map (
            O => \N__49638\,
            I => \N__49530\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__49631\,
            I => \N__49527\
        );

    \I__11696\ : InMux
    port map (
            O => \N__49630\,
            I => \N__49524\
        );

    \I__11695\ : CascadeMux
    port map (
            O => \N__49629\,
            I => \N__49518\
        );

    \I__11694\ : InMux
    port map (
            O => \N__49628\,
            I => \N__49515\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49512\
        );

    \I__11692\ : InMux
    port map (
            O => \N__49626\,
            I => \N__49509\
        );

    \I__11691\ : Span4Mux_h
    port map (
            O => \N__49623\,
            I => \N__49506\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__49620\,
            I => \N__49497\
        );

    \I__11689\ : Span4Mux_h
    port map (
            O => \N__49617\,
            I => \N__49497\
        );

    \I__11688\ : Span4Mux_v
    port map (
            O => \N__49614\,
            I => \N__49497\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__49605\,
            I => \N__49497\
        );

    \I__11686\ : Span4Mux_v
    port map (
            O => \N__49602\,
            I => \N__49492\
        );

    \I__11685\ : Span4Mux_v
    port map (
            O => \N__49599\,
            I => \N__49492\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49596\,
            I => \N__49489\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49595\,
            I => \N__49482\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49594\,
            I => \N__49482\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49482\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49592\,
            I => \N__49473\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49591\,
            I => \N__49473\
        );

    \I__11678\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49473\
        );

    \I__11677\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49473\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__49576\,
            I => \N__49462\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__49569\,
            I => \N__49462\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__49562\,
            I => \N__49462\
        );

    \I__11673\ : Span4Mux_v
    port map (
            O => \N__49555\,
            I => \N__49462\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__49548\,
            I => \N__49462\
        );

    \I__11671\ : Span4Mux_v
    port map (
            O => \N__49539\,
            I => \N__49457\
        );

    \I__11670\ : Span4Mux_v
    port map (
            O => \N__49536\,
            I => \N__49457\
        );

    \I__11669\ : Span4Mux_h
    port map (
            O => \N__49533\,
            I => \N__49450\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__49530\,
            I => \N__49450\
        );

    \I__11667\ : Span4Mux_h
    port map (
            O => \N__49527\,
            I => \N__49450\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__49524\,
            I => \N__49445\
        );

    \I__11665\ : InMux
    port map (
            O => \N__49523\,
            I => \N__49436\
        );

    \I__11664\ : InMux
    port map (
            O => \N__49522\,
            I => \N__49436\
        );

    \I__11663\ : InMux
    port map (
            O => \N__49521\,
            I => \N__49436\
        );

    \I__11662\ : InMux
    port map (
            O => \N__49518\,
            I => \N__49436\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__49515\,
            I => \N__49433\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__49512\,
            I => \N__49428\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__49509\,
            I => \N__49428\
        );

    \I__11658\ : Span4Mux_h
    port map (
            O => \N__49506\,
            I => \N__49423\
        );

    \I__11657\ : Span4Mux_v
    port map (
            O => \N__49497\,
            I => \N__49423\
        );

    \I__11656\ : Span4Mux_v
    port map (
            O => \N__49492\,
            I => \N__49418\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__49489\,
            I => \N__49418\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__49482\,
            I => \N__49407\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49407\
        );

    \I__11652\ : Span4Mux_h
    port map (
            O => \N__49462\,
            I => \N__49407\
        );

    \I__11651\ : Span4Mux_h
    port map (
            O => \N__49457\,
            I => \N__49407\
        );

    \I__11650\ : Span4Mux_h
    port map (
            O => \N__49450\,
            I => \N__49407\
        );

    \I__11649\ : InMux
    port map (
            O => \N__49449\,
            I => \N__49404\
        );

    \I__11648\ : InMux
    port map (
            O => \N__49448\,
            I => \N__49401\
        );

    \I__11647\ : Sp12to4
    port map (
            O => \N__49445\,
            I => \N__49396\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__49436\,
            I => \N__49396\
        );

    \I__11645\ : Span4Mux_h
    port map (
            O => \N__49433\,
            I => \N__49389\
        );

    \I__11644\ : Span4Mux_v
    port map (
            O => \N__49428\,
            I => \N__49389\
        );

    \I__11643\ : Span4Mux_v
    port map (
            O => \N__49423\,
            I => \N__49389\
        );

    \I__11642\ : Span4Mux_h
    port map (
            O => \N__49418\,
            I => \N__49384\
        );

    \I__11641\ : Span4Mux_v
    port map (
            O => \N__49407\,
            I => \N__49384\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__49404\,
            I => n9321
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__49401\,
            I => n9321
        );

    \I__11638\ : Odrv12
    port map (
            O => \N__49396\,
            I => n9321
        );

    \I__11637\ : Odrv4
    port map (
            O => \N__49389\,
            I => n9321
        );

    \I__11636\ : Odrv4
    port map (
            O => \N__49384\,
            I => n9321
        );

    \I__11635\ : InMux
    port map (
            O => \N__49373\,
            I => \N__49363\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49360\
        );

    \I__11633\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49345\
        );

    \I__11632\ : InMux
    port map (
            O => \N__49370\,
            I => \N__49345\
        );

    \I__11631\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49345\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49345\
        );

    \I__11629\ : InMux
    port map (
            O => \N__49367\,
            I => \N__49345\
        );

    \I__11628\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49339\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__49363\,
            I => \N__49336\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__49360\,
            I => \N__49333\
        );

    \I__11625\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49326\
        );

    \I__11624\ : InMux
    port map (
            O => \N__49358\,
            I => \N__49326\
        );

    \I__11623\ : InMux
    port map (
            O => \N__49357\,
            I => \N__49326\
        );

    \I__11622\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49323\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__49345\,
            I => \N__49320\
        );

    \I__11620\ : InMux
    port map (
            O => \N__49344\,
            I => \N__49317\
        );

    \I__11619\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49312\
        );

    \I__11618\ : InMux
    port map (
            O => \N__49342\,
            I => \N__49312\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__49339\,
            I => \N__49309\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__49336\,
            I => \N__49306\
        );

    \I__11615\ : Span4Mux_v
    port map (
            O => \N__49333\,
            I => \N__49303\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__49326\,
            I => \N__49296\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__49323\,
            I => \N__49296\
        );

    \I__11612\ : Span4Mux_h
    port map (
            O => \N__49320\,
            I => \N__49296\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__49317\,
            I => n12441
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__49312\,
            I => n12441
        );

    \I__11609\ : Odrv4
    port map (
            O => \N__49309\,
            I => n12441
        );

    \I__11608\ : Odrv4
    port map (
            O => \N__49306\,
            I => n12441
        );

    \I__11607\ : Odrv4
    port map (
            O => \N__49303\,
            I => n12441
        );

    \I__11606\ : Odrv4
    port map (
            O => \N__49296\,
            I => n12441
        );

    \I__11605\ : InMux
    port map (
            O => \N__49283\,
            I => \N__49279\
        );

    \I__11604\ : InMux
    port map (
            O => \N__49282\,
            I => \N__49276\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__49279\,
            I => \N__49272\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__49276\,
            I => \N__49269\
        );

    \I__11601\ : InMux
    port map (
            O => \N__49275\,
            I => \N__49266\
        );

    \I__11600\ : Span4Mux_h
    port map (
            O => \N__49272\,
            I => \N__49263\
        );

    \I__11599\ : Span4Mux_h
    port map (
            O => \N__49269\,
            I => \N__49260\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__49266\,
            I => \acadc_skipCount_4\
        );

    \I__11597\ : Odrv4
    port map (
            O => \N__49263\,
            I => \acadc_skipCount_4\
        );

    \I__11596\ : Odrv4
    port map (
            O => \N__49260\,
            I => \acadc_skipCount_4\
        );

    \I__11595\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49250\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__49250\,
            I => \N__49246\
        );

    \I__11593\ : CascadeMux
    port map (
            O => \N__49249\,
            I => \N__49243\
        );

    \I__11592\ : Span4Mux_h
    port map (
            O => \N__49246\,
            I => \N__49240\
        );

    \I__11591\ : InMux
    port map (
            O => \N__49243\,
            I => \N__49237\
        );

    \I__11590\ : Span4Mux_v
    port map (
            O => \N__49240\,
            I => \N__49234\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__49237\,
            I => data_idxvec_7
        );

    \I__11588\ : Odrv4
    port map (
            O => \N__49234\,
            I => data_idxvec_7
        );

    \I__11587\ : InMux
    port map (
            O => \N__49229\,
            I => \N__49226\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__49226\,
            I => \N__49221\
        );

    \I__11585\ : InMux
    port map (
            O => \N__49225\,
            I => \N__49218\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49224\,
            I => \N__49215\
        );

    \I__11583\ : Span4Mux_h
    port map (
            O => \N__49221\,
            I => \N__49212\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__49218\,
            I => data_cntvec_7
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__49215\,
            I => data_cntvec_7
        );

    \I__11580\ : Odrv4
    port map (
            O => \N__49212\,
            I => data_cntvec_7
        );

    \I__11579\ : InMux
    port map (
            O => \N__49205\,
            I => \N__49202\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__49202\,
            I => \N__49199\
        );

    \I__11577\ : Span4Mux_v
    port map (
            O => \N__49199\,
            I => \N__49196\
        );

    \I__11576\ : Odrv4
    port map (
            O => \N__49196\,
            I => buf_data_iac_15
        );

    \I__11575\ : CascadeMux
    port map (
            O => \N__49193\,
            I => \n26_adj_1500_cascade_\
        );

    \I__11574\ : CascadeMux
    port map (
            O => \N__49190\,
            I => \n20810_cascade_\
        );

    \I__11573\ : InMux
    port map (
            O => \N__49187\,
            I => \N__49184\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__49184\,
            I => n22058
        );

    \I__11571\ : CascadeMux
    port map (
            O => \N__49181\,
            I => \N__49177\
        );

    \I__11570\ : InMux
    port map (
            O => \N__49180\,
            I => \N__49173\
        );

    \I__11569\ : InMux
    port map (
            O => \N__49177\,
            I => \N__49170\
        );

    \I__11568\ : InMux
    port map (
            O => \N__49176\,
            I => \N__49167\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__49173\,
            I => \N__49162\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__49170\,
            I => \N__49162\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__49167\,
            I => \acadc_skipCount_7\
        );

    \I__11564\ : Odrv12
    port map (
            O => \N__49162\,
            I => \acadc_skipCount_7\
        );

    \I__11563\ : CascadeMux
    port map (
            O => \N__49157\,
            I => \N__49154\
        );

    \I__11562\ : InMux
    port map (
            O => \N__49154\,
            I => \N__49149\
        );

    \I__11561\ : InMux
    port map (
            O => \N__49153\,
            I => \N__49146\
        );

    \I__11560\ : InMux
    port map (
            O => \N__49152\,
            I => \N__49143\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__49149\,
            I => \N__49140\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__49146\,
            I => req_data_cnt_7
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__49143\,
            I => req_data_cnt_7
        );

    \I__11556\ : Odrv4
    port map (
            O => \N__49140\,
            I => req_data_cnt_7
        );

    \I__11555\ : InMux
    port map (
            O => \N__49133\,
            I => \N__49130\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__49130\,
            I => n20809
        );

    \I__11553\ : CascadeMux
    port map (
            O => \N__49127\,
            I => \N__49095\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49092\
        );

    \I__11551\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49089\
        );

    \I__11550\ : InMux
    port map (
            O => \N__49124\,
            I => \N__49086\
        );

    \I__11549\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49079\
        );

    \I__11548\ : InMux
    port map (
            O => \N__49122\,
            I => \N__49079\
        );

    \I__11547\ : InMux
    port map (
            O => \N__49121\,
            I => \N__49079\
        );

    \I__11546\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49069\
        );

    \I__11545\ : InMux
    port map (
            O => \N__49119\,
            I => \N__49069\
        );

    \I__11544\ : InMux
    port map (
            O => \N__49118\,
            I => \N__49066\
        );

    \I__11543\ : InMux
    port map (
            O => \N__49117\,
            I => \N__49063\
        );

    \I__11542\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49060\
        );

    \I__11541\ : InMux
    port map (
            O => \N__49115\,
            I => \N__49046\
        );

    \I__11540\ : InMux
    port map (
            O => \N__49114\,
            I => \N__49039\
        );

    \I__11539\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49039\
        );

    \I__11538\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49039\
        );

    \I__11537\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49030\
        );

    \I__11536\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49030\
        );

    \I__11535\ : InMux
    port map (
            O => \N__49109\,
            I => \N__49030\
        );

    \I__11534\ : InMux
    port map (
            O => \N__49108\,
            I => \N__49030\
        );

    \I__11533\ : InMux
    port map (
            O => \N__49107\,
            I => \N__49021\
        );

    \I__11532\ : InMux
    port map (
            O => \N__49106\,
            I => \N__49021\
        );

    \I__11531\ : InMux
    port map (
            O => \N__49105\,
            I => \N__49021\
        );

    \I__11530\ : InMux
    port map (
            O => \N__49104\,
            I => \N__49021\
        );

    \I__11529\ : InMux
    port map (
            O => \N__49103\,
            I => \N__49014\
        );

    \I__11528\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49014\
        );

    \I__11527\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49014\
        );

    \I__11526\ : InMux
    port map (
            O => \N__49100\,
            I => \N__49007\
        );

    \I__11525\ : InMux
    port map (
            O => \N__49099\,
            I => \N__49004\
        );

    \I__11524\ : InMux
    port map (
            O => \N__49098\,
            I => \N__49000\
        );

    \I__11523\ : InMux
    port map (
            O => \N__49095\,
            I => \N__48994\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__49092\,
            I => \N__48991\
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__49089\,
            I => \N__48984\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__49086\,
            I => \N__48984\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__49079\,
            I => \N__48984\
        );

    \I__11518\ : InMux
    port map (
            O => \N__49078\,
            I => \N__48977\
        );

    \I__11517\ : InMux
    port map (
            O => \N__49077\,
            I => \N__48977\
        );

    \I__11516\ : InMux
    port map (
            O => \N__49076\,
            I => \N__48977\
        );

    \I__11515\ : InMux
    port map (
            O => \N__49075\,
            I => \N__48974\
        );

    \I__11514\ : InMux
    port map (
            O => \N__49074\,
            I => \N__48971\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__49069\,
            I => \N__48966\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__49066\,
            I => \N__48966\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__49063\,
            I => \N__48961\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__48961\
        );

    \I__11509\ : InMux
    port map (
            O => \N__49059\,
            I => \N__48958\
        );

    \I__11508\ : InMux
    port map (
            O => \N__49058\,
            I => \N__48955\
        );

    \I__11507\ : InMux
    port map (
            O => \N__49057\,
            I => \N__48946\
        );

    \I__11506\ : InMux
    port map (
            O => \N__49056\,
            I => \N__48946\
        );

    \I__11505\ : InMux
    port map (
            O => \N__49055\,
            I => \N__48941\
        );

    \I__11504\ : InMux
    port map (
            O => \N__49054\,
            I => \N__48941\
        );

    \I__11503\ : InMux
    port map (
            O => \N__49053\,
            I => \N__48938\
        );

    \I__11502\ : InMux
    port map (
            O => \N__49052\,
            I => \N__48935\
        );

    \I__11501\ : InMux
    port map (
            O => \N__49051\,
            I => \N__48928\
        );

    \I__11500\ : InMux
    port map (
            O => \N__49050\,
            I => \N__48928\
        );

    \I__11499\ : InMux
    port map (
            O => \N__49049\,
            I => \N__48928\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__49046\,
            I => \N__48919\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__49039\,
            I => \N__48919\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__49030\,
            I => \N__48919\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48919\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__49014\,
            I => \N__48916\
        );

    \I__11493\ : InMux
    port map (
            O => \N__49013\,
            I => \N__48911\
        );

    \I__11492\ : InMux
    port map (
            O => \N__49012\,
            I => \N__48911\
        );

    \I__11491\ : InMux
    port map (
            O => \N__49011\,
            I => \N__48906\
        );

    \I__11490\ : InMux
    port map (
            O => \N__49010\,
            I => \N__48906\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__49007\,
            I => \N__48903\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48900\
        );

    \I__11487\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48897\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48894\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48887\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48887\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48997\,
            I => \N__48887\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__48994\,
            I => \N__48880\
        );

    \I__11481\ : Span4Mux_v
    port map (
            O => \N__48991\,
            I => \N__48880\
        );

    \I__11480\ : Span4Mux_v
    port map (
            O => \N__48984\,
            I => \N__48880\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__48977\,
            I => \N__48877\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__48974\,
            I => \N__48870\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48971\,
            I => \N__48865\
        );

    \I__11476\ : Span4Mux_v
    port map (
            O => \N__48966\,
            I => \N__48865\
        );

    \I__11475\ : Span4Mux_v
    port map (
            O => \N__48961\,
            I => \N__48860\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__48958\,
            I => \N__48860\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__48955\,
            I => \N__48857\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48954\,
            I => \N__48853\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48953\,
            I => \N__48846\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48952\,
            I => \N__48846\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48951\,
            I => \N__48846\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__48946\,
            I => \N__48841\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__48941\,
            I => \N__48841\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48938\,
            I => \N__48838\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48935\,
            I => \N__48835\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__48928\,
            I => \N__48826\
        );

    \I__11463\ : Span4Mux_v
    port map (
            O => \N__48919\,
            I => \N__48826\
        );

    \I__11462\ : Span4Mux_h
    port map (
            O => \N__48916\,
            I => \N__48826\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__48911\,
            I => \N__48826\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__48906\,
            I => \N__48817\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__48903\,
            I => \N__48817\
        );

    \I__11458\ : Span4Mux_h
    port map (
            O => \N__48900\,
            I => \N__48817\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__48897\,
            I => \N__48817\
        );

    \I__11456\ : Span4Mux_v
    port map (
            O => \N__48894\,
            I => \N__48810\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__48887\,
            I => \N__48810\
        );

    \I__11454\ : Span4Mux_h
    port map (
            O => \N__48880\,
            I => \N__48807\
        );

    \I__11453\ : Span12Mux_h
    port map (
            O => \N__48877\,
            I => \N__48804\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48795\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48875\,
            I => \N__48795\
        );

    \I__11450\ : InMux
    port map (
            O => \N__48874\,
            I => \N__48795\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48873\,
            I => \N__48795\
        );

    \I__11448\ : Span4Mux_v
    port map (
            O => \N__48870\,
            I => \N__48786\
        );

    \I__11447\ : Span4Mux_v
    port map (
            O => \N__48865\,
            I => \N__48786\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__48860\,
            I => \N__48786\
        );

    \I__11445\ : Span4Mux_v
    port map (
            O => \N__48857\,
            I => \N__48786\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48783\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48853\,
            I => \N__48776\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__48846\,
            I => \N__48776\
        );

    \I__11441\ : Span12Mux_v
    port map (
            O => \N__48841\,
            I => \N__48776\
        );

    \I__11440\ : Span4Mux_h
    port map (
            O => \N__48838\,
            I => \N__48767\
        );

    \I__11439\ : Span4Mux_v
    port map (
            O => \N__48835\,
            I => \N__48767\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__48826\,
            I => \N__48767\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__48817\,
            I => \N__48767\
        );

    \I__11436\ : InMux
    port map (
            O => \N__48816\,
            I => \N__48762\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48762\
        );

    \I__11434\ : Odrv4
    port map (
            O => \N__48810\,
            I => comm_cmd_2
        );

    \I__11433\ : Odrv4
    port map (
            O => \N__48807\,
            I => comm_cmd_2
        );

    \I__11432\ : Odrv12
    port map (
            O => \N__48804\,
            I => comm_cmd_2
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__48795\,
            I => comm_cmd_2
        );

    \I__11430\ : Odrv4
    port map (
            O => \N__48786\,
            I => comm_cmd_2
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__48783\,
            I => comm_cmd_2
        );

    \I__11428\ : Odrv12
    port map (
            O => \N__48776\,
            I => comm_cmd_2
        );

    \I__11427\ : Odrv4
    port map (
            O => \N__48767\,
            I => comm_cmd_2
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48762\,
            I => comm_cmd_2
        );

    \I__11425\ : CascadeMux
    port map (
            O => \N__48743\,
            I => \N__48731\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48724\
        );

    \I__11423\ : CascadeMux
    port map (
            O => \N__48741\,
            I => \N__48720\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48740\,
            I => \N__48715\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48709\
        );

    \I__11420\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48709\
        );

    \I__11419\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48704\
        );

    \I__11418\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48704\
        );

    \I__11417\ : InMux
    port map (
            O => \N__48735\,
            I => \N__48697\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48734\,
            I => \N__48692\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48731\,
            I => \N__48692\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48730\,
            I => \N__48689\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48729\,
            I => \N__48682\
        );

    \I__11412\ : CascadeMux
    port map (
            O => \N__48728\,
            I => \N__48678\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48727\,
            I => \N__48673\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__48724\,
            I => \N__48670\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48723\,
            I => \N__48665\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48662\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48719\,
            I => \N__48659\
        );

    \I__11406\ : CascadeMux
    port map (
            O => \N__48718\,
            I => \N__48656\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48715\,
            I => \N__48653\
        );

    \I__11404\ : InMux
    port map (
            O => \N__48714\,
            I => \N__48650\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__48709\,
            I => \N__48645\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__48704\,
            I => \N__48645\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48703\,
            I => \N__48642\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48702\,
            I => \N__48639\
        );

    \I__11399\ : InMux
    port map (
            O => \N__48701\,
            I => \N__48636\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48633\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48697\,
            I => \N__48626\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__48692\,
            I => \N__48626\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48689\,
            I => \N__48626\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48688\,
            I => \N__48621\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48687\,
            I => \N__48621\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48686\,
            I => \N__48614\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48614\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48611\
        );

    \I__11389\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48608\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48678\,
            I => \N__48602\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48677\,
            I => \N__48602\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48676\,
            I => \N__48599\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__48673\,
            I => \N__48594\
        );

    \I__11384\ : Span4Mux_v
    port map (
            O => \N__48670\,
            I => \N__48591\
        );

    \I__11383\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48588\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48585\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__48665\,
            I => \N__48578\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48578\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48659\,
            I => \N__48578\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48656\,
            I => \N__48575\
        );

    \I__11377\ : Span4Mux_h
    port map (
            O => \N__48653\,
            I => \N__48569\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__48650\,
            I => \N__48569\
        );

    \I__11375\ : Span4Mux_h
    port map (
            O => \N__48645\,
            I => \N__48564\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__48642\,
            I => \N__48564\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48639\,
            I => \N__48553\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48636\,
            I => \N__48553\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__48633\,
            I => \N__48553\
        );

    \I__11370\ : Span4Mux_v
    port map (
            O => \N__48626\,
            I => \N__48553\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__48621\,
            I => \N__48553\
        );

    \I__11368\ : CascadeMux
    port map (
            O => \N__48620\,
            I => \N__48550\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48619\,
            I => \N__48547\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__48614\,
            I => \N__48544\
        );

    \I__11365\ : Span4Mux_v
    port map (
            O => \N__48611\,
            I => \N__48539\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__48608\,
            I => \N__48539\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48607\,
            I => \N__48533\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__48602\,
            I => \N__48528\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__48599\,
            I => \N__48528\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48598\,
            I => \N__48523\
        );

    \I__11359\ : InMux
    port map (
            O => \N__48597\,
            I => \N__48523\
        );

    \I__11358\ : Span4Mux_h
    port map (
            O => \N__48594\,
            I => \N__48518\
        );

    \I__11357\ : Span4Mux_v
    port map (
            O => \N__48591\,
            I => \N__48518\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__48588\,
            I => \N__48515\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__48585\,
            I => \N__48510\
        );

    \I__11354\ : Span4Mux_h
    port map (
            O => \N__48578\,
            I => \N__48510\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48575\,
            I => \N__48507\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48574\,
            I => \N__48504\
        );

    \I__11351\ : Span4Mux_v
    port map (
            O => \N__48569\,
            I => \N__48496\
        );

    \I__11350\ : Span4Mux_v
    port map (
            O => \N__48564\,
            I => \N__48496\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__48553\,
            I => \N__48496\
        );

    \I__11348\ : InMux
    port map (
            O => \N__48550\,
            I => \N__48493\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__48547\,
            I => \N__48488\
        );

    \I__11346\ : Span4Mux_v
    port map (
            O => \N__48544\,
            I => \N__48488\
        );

    \I__11345\ : Span4Mux_h
    port map (
            O => \N__48539\,
            I => \N__48485\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48482\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48477\
        );

    \I__11342\ : InMux
    port map (
            O => \N__48536\,
            I => \N__48477\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__48533\,
            I => \N__48468\
        );

    \I__11340\ : Span12Mux_v
    port map (
            O => \N__48528\,
            I => \N__48468\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__48523\,
            I => \N__48468\
        );

    \I__11338\ : Sp12to4
    port map (
            O => \N__48518\,
            I => \N__48468\
        );

    \I__11337\ : Sp12to4
    port map (
            O => \N__48515\,
            I => \N__48465\
        );

    \I__11336\ : Span4Mux_v
    port map (
            O => \N__48510\,
            I => \N__48460\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__48507\,
            I => \N__48460\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__48504\,
            I => \N__48457\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48503\,
            I => \N__48454\
        );

    \I__11332\ : Span4Mux_h
    port map (
            O => \N__48496\,
            I => \N__48451\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__48493\,
            I => \N__48440\
        );

    \I__11330\ : Span4Mux_h
    port map (
            O => \N__48488\,
            I => \N__48440\
        );

    \I__11329\ : Span4Mux_v
    port map (
            O => \N__48485\,
            I => \N__48440\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__48482\,
            I => \N__48440\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__48477\,
            I => \N__48440\
        );

    \I__11326\ : Odrv12
    port map (
            O => \N__48468\,
            I => comm_cmd_3
        );

    \I__11325\ : Odrv12
    port map (
            O => \N__48465\,
            I => comm_cmd_3
        );

    \I__11324\ : Odrv4
    port map (
            O => \N__48460\,
            I => comm_cmd_3
        );

    \I__11323\ : Odrv12
    port map (
            O => \N__48457\,
            I => comm_cmd_3
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__48454\,
            I => comm_cmd_3
        );

    \I__11321\ : Odrv4
    port map (
            O => \N__48451\,
            I => comm_cmd_3
        );

    \I__11320\ : Odrv4
    port map (
            O => \N__48440\,
            I => comm_cmd_3
        );

    \I__11319\ : CascadeMux
    port map (
            O => \N__48425\,
            I => \N__48420\
        );

    \I__11318\ : CascadeMux
    port map (
            O => \N__48424\,
            I => \N__48411\
        );

    \I__11317\ : CascadeMux
    port map (
            O => \N__48423\,
            I => \N__48405\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48402\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48419\,
            I => \N__48399\
        );

    \I__11314\ : InMux
    port map (
            O => \N__48418\,
            I => \N__48395\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48417\,
            I => \N__48388\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48388\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48415\,
            I => \N__48388\
        );

    \I__11310\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48385\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48381\
        );

    \I__11308\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48378\
        );

    \I__11307\ : CascadeMux
    port map (
            O => \N__48409\,
            I => \N__48366\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48408\,
            I => \N__48354\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48405\,
            I => \N__48354\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48402\,
            I => \N__48351\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__48399\,
            I => \N__48348\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48398\,
            I => \N__48345\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__48395\,
            I => \N__48328\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48388\,
            I => \N__48328\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__48385\,
            I => \N__48328\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48325\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48322\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48319\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48305\
        );

    \I__11294\ : InMux
    port map (
            O => \N__48376\,
            I => \N__48300\
        );

    \I__11293\ : InMux
    port map (
            O => \N__48375\,
            I => \N__48300\
        );

    \I__11292\ : InMux
    port map (
            O => \N__48374\,
            I => \N__48289\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48286\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48278\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48371\,
            I => \N__48278\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48370\,
            I => \N__48278\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48369\,
            I => \N__48273\
        );

    \I__11286\ : InMux
    port map (
            O => \N__48366\,
            I => \N__48273\
        );

    \I__11285\ : CascadeMux
    port map (
            O => \N__48365\,
            I => \N__48270\
        );

    \I__11284\ : CascadeMux
    port map (
            O => \N__48364\,
            I => \N__48267\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48259\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48362\,
            I => \N__48259\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48361\,
            I => \N__48259\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48360\,
            I => \N__48256\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48359\,
            I => \N__48253\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__48354\,
            I => \N__48248\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__48351\,
            I => \N__48248\
        );

    \I__11276\ : Span4Mux_v
    port map (
            O => \N__48348\,
            I => \N__48243\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__48345\,
            I => \N__48243\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48344\,
            I => \N__48236\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48343\,
            I => \N__48236\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48236\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48233\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48229\
        );

    \I__11269\ : InMux
    port map (
            O => \N__48339\,
            I => \N__48223\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48223\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48337\,
            I => \N__48218\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48336\,
            I => \N__48218\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48335\,
            I => \N__48212\
        );

    \I__11264\ : Span4Mux_v
    port map (
            O => \N__48328\,
            I => \N__48203\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__48325\,
            I => \N__48203\
        );

    \I__11262\ : Span4Mux_h
    port map (
            O => \N__48322\,
            I => \N__48203\
        );

    \I__11261\ : Span4Mux_h
    port map (
            O => \N__48319\,
            I => \N__48203\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48196\
        );

    \I__11259\ : InMux
    port map (
            O => \N__48317\,
            I => \N__48196\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48316\,
            I => \N__48196\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48191\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48188\
        );

    \I__11255\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48185\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48312\,
            I => \N__48180\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48311\,
            I => \N__48180\
        );

    \I__11252\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48177\
        );

    \I__11251\ : InMux
    port map (
            O => \N__48309\,
            I => \N__48172\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48172\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48305\,
            I => \N__48167\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__48300\,
            I => \N__48164\
        );

    \I__11247\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48161\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48154\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48297\,
            I => \N__48154\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48296\,
            I => \N__48154\
        );

    \I__11243\ : InMux
    port map (
            O => \N__48295\,
            I => \N__48148\
        );

    \I__11242\ : InMux
    port map (
            O => \N__48294\,
            I => \N__48141\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48141\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48141\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__48289\,
            I => \N__48136\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48286\,
            I => \N__48136\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48133\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48278\,
            I => \N__48128\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__48273\,
            I => \N__48128\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48270\,
            I => \N__48123\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48123\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48120\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48117\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__48256\,
            I => \N__48114\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__48253\,
            I => \N__48111\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__48248\,
            I => \N__48102\
        );

    \I__11227\ : Span4Mux_v
    port map (
            O => \N__48243\,
            I => \N__48102\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__48236\,
            I => \N__48102\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48233\,
            I => \N__48102\
        );

    \I__11224\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48099\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__48229\,
            I => \N__48095\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48091\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48085\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48218\,
            I => \N__48085\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48078\
        );

    \I__11218\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48078\
        );

    \I__11217\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48078\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__48212\,
            I => \N__48073\
        );

    \I__11215\ : Span4Mux_h
    port map (
            O => \N__48203\,
            I => \N__48073\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48196\,
            I => \N__48070\
        );

    \I__11213\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48065\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48194\,
            I => \N__48065\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__48191\,
            I => \N__48054\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__48188\,
            I => \N__48054\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__48185\,
            I => \N__48054\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__48180\,
            I => \N__48054\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48177\,
            I => \N__48054\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48172\,
            I => \N__48051\
        );

    \I__11205\ : InMux
    port map (
            O => \N__48171\,
            I => \N__48046\
        );

    \I__11204\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48046\
        );

    \I__11203\ : Span4Mux_v
    port map (
            O => \N__48167\,
            I => \N__48037\
        );

    \I__11202\ : Span4Mux_h
    port map (
            O => \N__48164\,
            I => \N__48037\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__48161\,
            I => \N__48037\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48037\
        );

    \I__11199\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48030\
        );

    \I__11198\ : InMux
    port map (
            O => \N__48152\,
            I => \N__48030\
        );

    \I__11197\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48030\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__48148\,
            I => \N__48027\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__48024\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__48136\,
            I => \N__48021\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__48133\,
            I => \N__48014\
        );

    \I__11192\ : Span4Mux_v
    port map (
            O => \N__48128\,
            I => \N__48014\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__48123\,
            I => \N__48014\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__48120\,
            I => \N__48011\
        );

    \I__11189\ : Span4Mux_h
    port map (
            O => \N__48117\,
            I => \N__48008\
        );

    \I__11188\ : Span4Mux_h
    port map (
            O => \N__48114\,
            I => \N__47999\
        );

    \I__11187\ : Span4Mux_h
    port map (
            O => \N__48111\,
            I => \N__47999\
        );

    \I__11186\ : Span4Mux_h
    port map (
            O => \N__48102\,
            I => \N__47999\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__47999\
        );

    \I__11184\ : InMux
    port map (
            O => \N__48098\,
            I => \N__47994\
        );

    \I__11183\ : Span4Mux_h
    port map (
            O => \N__48095\,
            I => \N__47991\
        );

    \I__11182\ : InMux
    port map (
            O => \N__48094\,
            I => \N__47988\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__48091\,
            I => \N__47985\
        );

    \I__11180\ : InMux
    port map (
            O => \N__48090\,
            I => \N__47982\
        );

    \I__11179\ : Span4Mux_h
    port map (
            O => \N__48085\,
            I => \N__47975\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__48078\,
            I => \N__47975\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__48073\,
            I => \N__47975\
        );

    \I__11176\ : Span4Mux_h
    port map (
            O => \N__48070\,
            I => \N__47970\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__48065\,
            I => \N__47970\
        );

    \I__11174\ : Span4Mux_v
    port map (
            O => \N__48054\,
            I => \N__47961\
        );

    \I__11173\ : Span4Mux_v
    port map (
            O => \N__48051\,
            I => \N__47961\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__48046\,
            I => \N__47961\
        );

    \I__11171\ : Span4Mux_v
    port map (
            O => \N__48037\,
            I => \N__47961\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__48030\,
            I => \N__47950\
        );

    \I__11169\ : Span4Mux_v
    port map (
            O => \N__48027\,
            I => \N__47950\
        );

    \I__11168\ : Span4Mux_v
    port map (
            O => \N__48024\,
            I => \N__47950\
        );

    \I__11167\ : Span4Mux_h
    port map (
            O => \N__48021\,
            I => \N__47950\
        );

    \I__11166\ : Span4Mux_v
    port map (
            O => \N__48014\,
            I => \N__47950\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__48011\,
            I => \N__47943\
        );

    \I__11164\ : Span4Mux_v
    port map (
            O => \N__48008\,
            I => \N__47943\
        );

    \I__11163\ : Span4Mux_v
    port map (
            O => \N__47999\,
            I => \N__47943\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47998\,
            I => \N__47938\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47938\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47994\,
            I => comm_cmd_1
        );

    \I__11159\ : Odrv4
    port map (
            O => \N__47991\,
            I => comm_cmd_1
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__47988\,
            I => comm_cmd_1
        );

    \I__11157\ : Odrv12
    port map (
            O => \N__47985\,
            I => comm_cmd_1
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__47982\,
            I => comm_cmd_1
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47975\,
            I => comm_cmd_1
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__47970\,
            I => comm_cmd_1
        );

    \I__11153\ : Odrv4
    port map (
            O => \N__47961\,
            I => comm_cmd_1
        );

    \I__11152\ : Odrv4
    port map (
            O => \N__47950\,
            I => comm_cmd_1
        );

    \I__11151\ : Odrv4
    port map (
            O => \N__47943\,
            I => comm_cmd_1
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__47938\,
            I => comm_cmd_1
        );

    \I__11149\ : CascadeMux
    port map (
            O => \N__47915\,
            I => \N__47912\
        );

    \I__11148\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47908\
        );

    \I__11147\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47905\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47908\,
            I => \N__47902\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__47905\,
            I => \N__47899\
        );

    \I__11144\ : Span4Mux_v
    port map (
            O => \N__47902\,
            I => \N__47894\
        );

    \I__11143\ : Span4Mux_h
    port map (
            O => \N__47899\,
            I => \N__47894\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__47894\,
            I => \N__47891\
        );

    \I__11141\ : Odrv4
    port map (
            O => \N__47891\,
            I => comm_length_1
        );

    \I__11140\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47884\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47881\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__47884\,
            I => comm_length_2
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__47881\,
            I => comm_length_2
        );

    \I__11136\ : CascadeMux
    port map (
            O => \N__47876\,
            I => \N__47873\
        );

    \I__11135\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47870\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__47870\,
            I => comm_length_0
        );

    \I__11133\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47863\
        );

    \I__11132\ : InMux
    port map (
            O => \N__47866\,
            I => \N__47860\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__47863\,
            I => \N__47857\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47860\,
            I => \N__47854\
        );

    \I__11129\ : Span4Mux_v
    port map (
            O => \N__47857\,
            I => \N__47851\
        );

    \I__11128\ : Span12Mux_v
    port map (
            O => \N__47854\,
            I => \N__47848\
        );

    \I__11127\ : Odrv4
    port map (
            O => \N__47851\,
            I => n4
        );

    \I__11126\ : Odrv12
    port map (
            O => \N__47848\,
            I => n4
        );

    \I__11125\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47838\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47835\
        );

    \I__11123\ : CascadeMux
    port map (
            O => \N__47841\,
            I => \N__47832\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__47838\,
            I => \N__47829\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47835\,
            I => \N__47826\
        );

    \I__11120\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47823\
        );

    \I__11119\ : Span4Mux_v
    port map (
            O => \N__47829\,
            I => \N__47818\
        );

    \I__11118\ : Span4Mux_h
    port map (
            O => \N__47826\,
            I => \N__47818\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__47823\,
            I => \N__47815\
        );

    \I__11116\ : Span4Mux_h
    port map (
            O => \N__47818\,
            I => \N__47812\
        );

    \I__11115\ : Span4Mux_h
    port map (
            O => \N__47815\,
            I => \N__47809\
        );

    \I__11114\ : Span4Mux_h
    port map (
            O => \N__47812\,
            I => \N__47806\
        );

    \I__11113\ : Span4Mux_v
    port map (
            O => \N__47809\,
            I => \N__47803\
        );

    \I__11112\ : Span4Mux_v
    port map (
            O => \N__47806\,
            I => \N__47800\
        );

    \I__11111\ : Odrv4
    port map (
            O => \N__47803\,
            I => n14_adj_1579
        );

    \I__11110\ : Odrv4
    port map (
            O => \N__47800\,
            I => n14_adj_1579
        );

    \I__11109\ : CascadeMux
    port map (
            O => \N__47795\,
            I => \N__47791\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47788\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47784\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47781\
        );

    \I__11105\ : CascadeMux
    port map (
            O => \N__47787\,
            I => \N__47778\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47784\,
            I => \N__47773\
        );

    \I__11103\ : Span4Mux_h
    port map (
            O => \N__47781\,
            I => \N__47773\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47770\
        );

    \I__11101\ : Odrv4
    port map (
            O => \N__47773\,
            I => \acadc_skipCount_15\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__47770\,
            I => \acadc_skipCount_15\
        );

    \I__11099\ : CascadeMux
    port map (
            O => \N__47765\,
            I => \N__47762\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47756\
        );

    \I__11096\ : Odrv12
    port map (
            O => \N__47756\,
            I => n23_adj_1527
        );

    \I__11095\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47749\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47752\,
            I => \N__47746\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__47749\,
            I => \N__47740\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47746\,
            I => \N__47740\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47737\
        );

    \I__11090\ : Odrv12
    port map (
            O => \N__47740\,
            I => data_cntvec_5
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__47737\,
            I => data_cntvec_5
        );

    \I__11088\ : InMux
    port map (
            O => \N__47732\,
            I => \N__47727\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47724\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47721\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47727\,
            I => \N__47718\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47715\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__47721\,
            I => data_cntvec_3
        );

    \I__11082\ : Odrv4
    port map (
            O => \N__47718\,
            I => data_cntvec_3
        );

    \I__11081\ : Odrv4
    port map (
            O => \N__47715\,
            I => data_cntvec_3
        );

    \I__11080\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47705\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47705\,
            I => \N__47702\
        );

    \I__11078\ : Span4Mux_h
    port map (
            O => \N__47702\,
            I => \N__47697\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47692\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47692\
        );

    \I__11075\ : Odrv4
    port map (
            O => \N__47697\,
            I => req_data_cnt_3
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47692\,
            I => req_data_cnt_3
        );

    \I__11073\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47684\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47684\,
            I => n20_adj_1596
        );

    \I__11071\ : CascadeMux
    port map (
            O => \N__47681\,
            I => \N__47677\
        );

    \I__11070\ : CascadeMux
    port map (
            O => \N__47680\,
            I => \N__47674\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47669\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47666\
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__47673\,
            I => \N__47663\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47660\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47657\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__47666\,
            I => \N__47653\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47663\,
            I => \N__47650\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__47660\,
            I => \N__47647\
        );

    \I__11061\ : Span4Mux_v
    port map (
            O => \N__47657\,
            I => \N__47644\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47656\,
            I => \N__47641\
        );

    \I__11059\ : Span4Mux_v
    port map (
            O => \N__47653\,
            I => \N__47634\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47634\
        );

    \I__11057\ : Span4Mux_h
    port map (
            O => \N__47647\,
            I => \N__47634\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__47644\,
            I => \N__47631\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47641\,
            I => \N__47627\
        );

    \I__11054\ : Span4Mux_h
    port map (
            O => \N__47634\,
            I => \N__47624\
        );

    \I__11053\ : Span4Mux_h
    port map (
            O => \N__47631\,
            I => \N__47621\
        );

    \I__11052\ : InMux
    port map (
            O => \N__47630\,
            I => \N__47618\
        );

    \I__11051\ : Span4Mux_v
    port map (
            O => \N__47627\,
            I => \N__47613\
        );

    \I__11050\ : Span4Mux_v
    port map (
            O => \N__47624\,
            I => \N__47613\
        );

    \I__11049\ : Odrv4
    port map (
            O => \N__47621\,
            I => comm_buf_1_7
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47618\,
            I => comm_buf_1_7
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__47613\,
            I => comm_buf_1_7
        );

    \I__11046\ : InMux
    port map (
            O => \N__47606\,
            I => \N__47603\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47603\,
            I => \N__47600\
        );

    \I__11044\ : Span12Mux_v
    port map (
            O => \N__47600\,
            I => \N__47597\
        );

    \I__11043\ : Odrv12
    port map (
            O => \N__47597\,
            I => n14_adj_1546
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__47594\,
            I => \n14_adj_1546_cascade_\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__47591\,
            I => \N__47588\
        );

    \I__11040\ : InMux
    port map (
            O => \N__47588\,
            I => \N__47584\
        );

    \I__11039\ : InMux
    port map (
            O => \N__47587\,
            I => \N__47581\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__47584\,
            I => \N__47576\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__47581\,
            I => \N__47576\
        );

    \I__11036\ : Span4Mux_v
    port map (
            O => \N__47576\,
            I => \N__47572\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47575\,
            I => \N__47569\
        );

    \I__11034\ : Span4Mux_h
    port map (
            O => \N__47572\,
            I => \N__47566\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__47569\,
            I => \N__47563\
        );

    \I__11032\ : Sp12to4
    port map (
            O => \N__47566\,
            I => \N__47560\
        );

    \I__11031\ : Odrv12
    port map (
            O => \N__47563\,
            I => n14_adj_1577
        );

    \I__11030\ : Odrv12
    port map (
            O => \N__47560\,
            I => n14_adj_1577
        );

    \I__11029\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47552\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__47552\,
            I => \N__47548\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47551\,
            I => \N__47544\
        );

    \I__11026\ : Span12Mux_h
    port map (
            O => \N__47548\,
            I => \N__47541\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47547\,
            I => \N__47538\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47544\,
            I => req_data_cnt_13
        );

    \I__11023\ : Odrv12
    port map (
            O => \N__47541\,
            I => req_data_cnt_13
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__47538\,
            I => req_data_cnt_13
        );

    \I__11021\ : InMux
    port map (
            O => \N__47531\,
            I => \N__47527\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47530\,
            I => \N__47523\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__47527\,
            I => \N__47520\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47526\,
            I => \N__47517\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__47523\,
            I => data_cntvec_9
        );

    \I__11016\ : Odrv4
    port map (
            O => \N__47520\,
            I => data_cntvec_9
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47517\,
            I => data_cntvec_9
        );

    \I__11014\ : InMux
    port map (
            O => \N__47510\,
            I => \N__47507\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47503\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47506\,
            I => \N__47499\
        );

    \I__11011\ : Span4Mux_h
    port map (
            O => \N__47503\,
            I => \N__47496\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47493\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__47499\,
            I => req_data_cnt_15
        );

    \I__11008\ : Odrv4
    port map (
            O => \N__47496\,
            I => req_data_cnt_15
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__47493\,
            I => req_data_cnt_15
        );

    \I__11006\ : CascadeMux
    port map (
            O => \N__47486\,
            I => \N__47482\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47485\,
            I => \N__47479\
        );

    \I__11004\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47476\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47479\,
            I => \N__47471\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__47476\,
            I => \N__47471\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__47471\,
            I => data_cntvec_15
        );

    \I__11000\ : InMux
    port map (
            O => \N__47468\,
            I => \N__47465\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__47465\,
            I => n24
        );

    \I__10998\ : InMux
    port map (
            O => \N__47462\,
            I => \N__47458\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47455\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47452\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__47455\,
            I => \N__47449\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__47452\,
            I => \N__47446\
        );

    \I__10993\ : Sp12to4
    port map (
            O => \N__47449\,
            I => \N__47443\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__47446\,
            I => \N__47440\
        );

    \I__10991\ : Span12Mux_v
    port map (
            O => \N__47443\,
            I => \N__47437\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__47440\,
            I => n14_adj_1574
        );

    \I__10989\ : Odrv12
    port map (
            O => \N__47437\,
            I => n14_adj_1574
        );

    \I__10988\ : InMux
    port map (
            O => \N__47432\,
            I => \N__47429\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__47429\,
            I => \N__47424\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47419\
        );

    \I__10985\ : InMux
    port map (
            O => \N__47427\,
            I => \N__47419\
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__47424\,
            I => req_data_cnt_9
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47419\,
            I => req_data_cnt_9
        );

    \I__10982\ : InMux
    port map (
            O => \N__47414\,
            I => \N__47406\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47406\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47401\
        );

    \I__10979\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47401\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47406\,
            I => \N__47398\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__47401\,
            I => \N__47392\
        );

    \I__10976\ : Span4Mux_h
    port map (
            O => \N__47398\,
            I => \N__47389\
        );

    \I__10975\ : InMux
    port map (
            O => \N__47397\,
            I => \N__47382\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47396\,
            I => \N__47382\
        );

    \I__10973\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47382\
        );

    \I__10972\ : Span4Mux_v
    port map (
            O => \N__47392\,
            I => \N__47372\
        );

    \I__10971\ : Span4Mux_h
    port map (
            O => \N__47389\,
            I => \N__47367\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__47382\,
            I => \N__47367\
        );

    \I__10969\ : InMux
    port map (
            O => \N__47381\,
            I => \N__47358\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47358\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47358\
        );

    \I__10966\ : InMux
    port map (
            O => \N__47378\,
            I => \N__47358\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47351\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47376\,
            I => \N__47351\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47375\,
            I => \N__47351\
        );

    \I__10962\ : Span4Mux_h
    port map (
            O => \N__47372\,
            I => \N__47347\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__47367\,
            I => \N__47344\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__47358\,
            I => \N__47339\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__47351\,
            I => \N__47339\
        );

    \I__10958\ : InMux
    port map (
            O => \N__47350\,
            I => \N__47336\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__47347\,
            I => n12467
        );

    \I__10956\ : Odrv4
    port map (
            O => \N__47344\,
            I => n12467
        );

    \I__10955\ : Odrv12
    port map (
            O => \N__47339\,
            I => n12467
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__47336\,
            I => n12467
        );

    \I__10953\ : CascadeMux
    port map (
            O => \N__47327\,
            I => \N__47323\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47326\,
            I => \N__47319\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47316\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47313\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47319\,
            I => \N__47310\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47316\,
            I => \N__47307\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__47313\,
            I => \N__47304\
        );

    \I__10946\ : Span4Mux_v
    port map (
            O => \N__47310\,
            I => \N__47301\
        );

    \I__10945\ : Span12Mux_v
    port map (
            O => \N__47307\,
            I => \N__47296\
        );

    \I__10944\ : Span12Mux_h
    port map (
            O => \N__47304\,
            I => \N__47296\
        );

    \I__10943\ : Odrv4
    port map (
            O => \N__47301\,
            I => n14_adj_1578
        );

    \I__10942\ : Odrv12
    port map (
            O => \N__47296\,
            I => n14_adj_1578
        );

    \I__10941\ : CascadeMux
    port map (
            O => \N__47291\,
            I => \N__47288\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47288\,
            I => \N__47285\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47285\,
            I => \N__47280\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__47284\,
            I => \N__47277\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47283\,
            I => \N__47274\
        );

    \I__10936\ : Span4Mux_v
    port map (
            O => \N__47280\,
            I => \N__47271\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47268\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47274\,
            I => \N__47263\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__47271\,
            I => \N__47263\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47268\,
            I => \N__47260\
        );

    \I__10931\ : Odrv4
    port map (
            O => \N__47263\,
            I => req_data_cnt_5
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__47260\,
            I => req_data_cnt_5
        );

    \I__10929\ : CascadeMux
    port map (
            O => \N__47255\,
            I => \n22211_cascade_\
        );

    \I__10928\ : CascadeMux
    port map (
            O => \N__47252\,
            I => \N__47249\
        );

    \I__10927\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47243\
        );

    \I__10926\ : CascadeMux
    port map (
            O => \N__47248\,
            I => \N__47238\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47235\
        );

    \I__10924\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47231\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__47243\,
            I => \N__47228\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47242\,
            I => \N__47225\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47222\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47238\,
            I => \N__47218\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__47235\,
            I => \N__47215\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47212\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47231\,
            I => \N__47209\
        );

    \I__10916\ : Span4Mux_v
    port map (
            O => \N__47228\,
            I => \N__47202\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__47225\,
            I => \N__47202\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__47222\,
            I => \N__47202\
        );

    \I__10913\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47199\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47218\,
            I => \N__47196\
        );

    \I__10911\ : Sp12to4
    port map (
            O => \N__47215\,
            I => \N__47191\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47191\
        );

    \I__10909\ : Span4Mux_v
    port map (
            O => \N__47209\,
            I => \N__47188\
        );

    \I__10908\ : Span4Mux_v
    port map (
            O => \N__47202\,
            I => \N__47185\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__47199\,
            I => \N__47182\
        );

    \I__10906\ : Span12Mux_h
    port map (
            O => \N__47196\,
            I => \N__47178\
        );

    \I__10905\ : Span12Mux_v
    port map (
            O => \N__47191\,
            I => \N__47175\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__47188\,
            I => \N__47170\
        );

    \I__10903\ : Span4Mux_v
    port map (
            O => \N__47185\,
            I => \N__47170\
        );

    \I__10902\ : Span4Mux_h
    port map (
            O => \N__47182\,
            I => \N__47167\
        );

    \I__10901\ : InMux
    port map (
            O => \N__47181\,
            I => \N__47164\
        );

    \I__10900\ : Odrv12
    port map (
            O => \N__47178\,
            I => comm_rx_buf_2
        );

    \I__10899\ : Odrv12
    port map (
            O => \N__47175\,
            I => comm_rx_buf_2
        );

    \I__10898\ : Odrv4
    port map (
            O => \N__47170\,
            I => comm_rx_buf_2
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__47167\,
            I => comm_rx_buf_2
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47164\,
            I => comm_rx_buf_2
        );

    \I__10895\ : CascadeMux
    port map (
            O => \N__47153\,
            I => \n30_adj_1518_cascade_\
        );

    \I__10894\ : CascadeMux
    port map (
            O => \N__47150\,
            I => \N__47147\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47144\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__47144\,
            I => \N__47140\
        );

    \I__10891\ : CascadeMux
    port map (
            O => \N__47143\,
            I => \N__47136\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__47140\,
            I => \N__47130\
        );

    \I__10889\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47127\
        );

    \I__10888\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47124\
        );

    \I__10887\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47121\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47118\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47115\
        );

    \I__10884\ : Span4Mux_h
    port map (
            O => \N__47130\,
            I => \N__47110\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__47127\,
            I => \N__47110\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__47124\,
            I => \N__47105\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__47121\,
            I => \N__47105\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__47118\,
            I => \N__47102\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47115\,
            I => \N__47099\
        );

    \I__10878\ : Span4Mux_v
    port map (
            O => \N__47110\,
            I => \N__47096\
        );

    \I__10877\ : Span12Mux_h
    port map (
            O => \N__47105\,
            I => \N__47093\
        );

    \I__10876\ : Span4Mux_h
    port map (
            O => \N__47102\,
            I => \N__47090\
        );

    \I__10875\ : Span4Mux_v
    port map (
            O => \N__47099\,
            I => \N__47087\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__47096\,
            I => \N__47084\
        );

    \I__10873\ : Odrv12
    port map (
            O => \N__47093\,
            I => comm_buf_1_2
        );

    \I__10872\ : Odrv4
    port map (
            O => \N__47090\,
            I => comm_buf_1_2
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__47087\,
            I => comm_buf_1_2
        );

    \I__10870\ : Odrv4
    port map (
            O => \N__47084\,
            I => comm_buf_1_2
        );

    \I__10869\ : CEMux
    port map (
            O => \N__47075\,
            I => \N__47072\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__47072\,
            I => \N__47065\
        );

    \I__10867\ : CEMux
    port map (
            O => \N__47071\,
            I => \N__47062\
        );

    \I__10866\ : CEMux
    port map (
            O => \N__47070\,
            I => \N__47058\
        );

    \I__10865\ : CEMux
    port map (
            O => \N__47069\,
            I => \N__47055\
        );

    \I__10864\ : CEMux
    port map (
            O => \N__47068\,
            I => \N__47050\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__47065\,
            I => \N__47045\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__47062\,
            I => \N__47045\
        );

    \I__10861\ : CEMux
    port map (
            O => \N__47061\,
            I => \N__47042\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__47058\,
            I => \N__47039\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47036\
        );

    \I__10858\ : CEMux
    port map (
            O => \N__47054\,
            I => \N__47033\
        );

    \I__10857\ : CEMux
    port map (
            O => \N__47053\,
            I => \N__47030\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__47050\,
            I => \N__47022\
        );

    \I__10855\ : Span4Mux_h
    port map (
            O => \N__47045\,
            I => \N__47022\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__47042\,
            I => \N__47022\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__47039\,
            I => \N__47015\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__47036\,
            I => \N__47015\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__47033\,
            I => \N__47015\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47012\
        );

    \I__10849\ : InMux
    port map (
            O => \N__47029\,
            I => \N__47009\
        );

    \I__10848\ : Odrv4
    port map (
            O => \N__47022\,
            I => n12047
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__47015\,
            I => n12047
        );

    \I__10846\ : Odrv12
    port map (
            O => \N__47012\,
            I => n12047
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__47009\,
            I => n12047
        );

    \I__10844\ : SRMux
    port map (
            O => \N__47000\,
            I => \N__46997\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46990\
        );

    \I__10842\ : SRMux
    port map (
            O => \N__46996\,
            I => \N__46986\
        );

    \I__10841\ : SRMux
    port map (
            O => \N__46995\,
            I => \N__46983\
        );

    \I__10840\ : SRMux
    port map (
            O => \N__46994\,
            I => \N__46980\
        );

    \I__10839\ : SRMux
    port map (
            O => \N__46993\,
            I => \N__46977\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__46990\,
            I => \N__46974\
        );

    \I__10837\ : SRMux
    port map (
            O => \N__46989\,
            I => \N__46971\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46986\,
            I => \N__46966\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__46983\,
            I => \N__46963\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46980\,
            I => \N__46960\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46957\
        );

    \I__10832\ : Span4Mux_h
    port map (
            O => \N__46974\,
            I => \N__46952\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__46971\,
            I => \N__46952\
        );

    \I__10830\ : SRMux
    port map (
            O => \N__46970\,
            I => \N__46949\
        );

    \I__10829\ : SRMux
    port map (
            O => \N__46969\,
            I => \N__46946\
        );

    \I__10828\ : Span4Mux_v
    port map (
            O => \N__46966\,
            I => \N__46941\
        );

    \I__10827\ : Span4Mux_v
    port map (
            O => \N__46963\,
            I => \N__46941\
        );

    \I__10826\ : Span4Mux_v
    port map (
            O => \N__46960\,
            I => \N__46936\
        );

    \I__10825\ : Span4Mux_h
    port map (
            O => \N__46957\,
            I => \N__46936\
        );

    \I__10824\ : Span4Mux_h
    port map (
            O => \N__46952\,
            I => \N__46933\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46949\,
            I => \N__46930\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46927\
        );

    \I__10821\ : Odrv4
    port map (
            O => \N__46941\,
            I => n14773
        );

    \I__10820\ : Odrv4
    port map (
            O => \N__46936\,
            I => n14773
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__46933\,
            I => n14773
        );

    \I__10818\ : Odrv12
    port map (
            O => \N__46930\,
            I => n14773
        );

    \I__10817\ : Odrv12
    port map (
            O => \N__46927\,
            I => n14773
        );

    \I__10816\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46913\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46913\,
            I => \N__46910\
        );

    \I__10814\ : Span4Mux_h
    port map (
            O => \N__46910\,
            I => \N__46907\
        );

    \I__10813\ : Span4Mux_h
    port map (
            O => \N__46907\,
            I => \N__46904\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__46904\,
            I => n19_adj_1516
        );

    \I__10811\ : CascadeMux
    port map (
            O => \N__46901\,
            I => \N__46898\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46895\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46892\
        );

    \I__10808\ : Span12Mux_h
    port map (
            O => \N__46892\,
            I => \N__46888\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46885\
        );

    \I__10806\ : Odrv12
    port map (
            O => \N__46888\,
            I => \buf_readRTD_2\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46885\,
            I => \buf_readRTD_2\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46877\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46877\,
            I => n21956
        );

    \I__10802\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46871\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46871\,
            I => \N__46867\
        );

    \I__10800\ : CascadeMux
    port map (
            O => \N__46870\,
            I => \N__46864\
        );

    \I__10799\ : Span4Mux_h
    port map (
            O => \N__46867\,
            I => \N__46861\
        );

    \I__10798\ : InMux
    port map (
            O => \N__46864\,
            I => \N__46858\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__46861\,
            I => \N__46855\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__46858\,
            I => data_idxvec_2
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__46855\,
            I => data_idxvec_2
        );

    \I__10794\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46846\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46842\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46839\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46845\,
            I => \N__46836\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46842\,
            I => \N__46833\
        );

    \I__10789\ : Span4Mux_h
    port map (
            O => \N__46839\,
            I => \N__46830\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46836\,
            I => data_cntvec_2
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__46833\,
            I => data_cntvec_2
        );

    \I__10786\ : Odrv4
    port map (
            O => \N__46830\,
            I => data_cntvec_2
        );

    \I__10785\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46820\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__46820\,
            I => n26_adj_1517
        );

    \I__10783\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46813\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46810\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46813\,
            I => \N__46807\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__46810\,
            I => \N__46804\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__46807\,
            I => \N__46799\
        );

    \I__10778\ : Span4Mux_v
    port map (
            O => \N__46804\,
            I => \N__46799\
        );

    \I__10777\ : Odrv4
    port map (
            O => \N__46799\,
            I => n14_adj_1550
        );

    \I__10776\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46792\
        );

    \I__10775\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46789\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__46792\,
            I => \N__46786\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__46789\,
            I => \N__46783\
        );

    \I__10772\ : Span4Mux_h
    port map (
            O => \N__46786\,
            I => \N__46780\
        );

    \I__10771\ : Span4Mux_h
    port map (
            O => \N__46783\,
            I => \N__46777\
        );

    \I__10770\ : Odrv4
    port map (
            O => \N__46780\,
            I => n14_adj_1544
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__46777\,
            I => n14_adj_1544
        );

    \I__10768\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46769\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__46769\,
            I => \N__46764\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46761\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46758\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__46764\,
            I => \N__46755\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46761\,
            I => \N__46752\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46758\,
            I => data_cntvec_1
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__46755\,
            I => data_cntvec_1
        );

    \I__10760\ : Odrv4
    port map (
            O => \N__46752\,
            I => data_cntvec_1
        );

    \I__10759\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46741\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46737\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__46741\,
            I => \N__46734\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46731\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__46737\,
            I => data_cntvec_4
        );

    \I__10754\ : Odrv4
    port map (
            O => \N__46734\,
            I => data_cntvec_4
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__46731\,
            I => data_cntvec_4
        );

    \I__10752\ : InMux
    port map (
            O => \N__46724\,
            I => \N__46720\
        );

    \I__10751\ : CascadeMux
    port map (
            O => \N__46723\,
            I => \N__46717\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46713\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46710\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46707\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__46713\,
            I => \N__46704\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__46710\,
            I => \N__46701\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__46707\,
            I => req_data_cnt_4
        );

    \I__10744\ : Odrv4
    port map (
            O => \N__46704\,
            I => req_data_cnt_4
        );

    \I__10743\ : Odrv4
    port map (
            O => \N__46701\,
            I => req_data_cnt_4
        );

    \I__10742\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46691\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46686\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46690\,
            I => \N__46681\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46681\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__46686\,
            I => req_data_cnt_1
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46681\,
            I => req_data_cnt_1
        );

    \I__10736\ : InMux
    port map (
            O => \N__46676\,
            I => \N__46673\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__46673\,
            I => n18
        );

    \I__10734\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46667\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46667\,
            I => \N__46663\
        );

    \I__10732\ : CascadeMux
    port map (
            O => \N__46666\,
            I => \N__46660\
        );

    \I__10731\ : Span12Mux_v
    port map (
            O => \N__46663\,
            I => \N__46657\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46654\
        );

    \I__10729\ : Odrv12
    port map (
            O => \N__46657\,
            I => buf_adcdata_vdc_13
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__46654\,
            I => buf_adcdata_vdc_13
        );

    \I__10727\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46646\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__46646\,
            I => \N__46643\
        );

    \I__10725\ : Span4Mux_v
    port map (
            O => \N__46643\,
            I => \N__46639\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46636\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__46639\,
            I => \N__46630\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46636\,
            I => \N__46630\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46635\,
            I => \N__46627\
        );

    \I__10720\ : Span4Mux_h
    port map (
            O => \N__46630\,
            I => \N__46624\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__46627\,
            I => buf_adcdata_vac_13
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__46624\,
            I => buf_adcdata_vac_13
        );

    \I__10717\ : InMux
    port map (
            O => \N__46619\,
            I => \N__46616\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46616\,
            I => n19_adj_1497
        );

    \I__10715\ : InMux
    port map (
            O => \N__46613\,
            I => \N__46610\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46606\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46609\,
            I => \N__46603\
        );

    \I__10712\ : Span4Mux_v
    port map (
            O => \N__46606\,
            I => \N__46600\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46597\
        );

    \I__10710\ : Sp12to4
    port map (
            O => \N__46600\,
            I => \N__46594\
        );

    \I__10709\ : Span4Mux_h
    port map (
            O => \N__46597\,
            I => \N__46591\
        );

    \I__10708\ : Odrv12
    port map (
            O => \N__46594\,
            I => n9
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__46591\,
            I => n9
        );

    \I__10706\ : InMux
    port map (
            O => \N__46586\,
            I => \N__46582\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46578\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__46582\,
            I => \N__46575\
        );

    \I__10703\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46572\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__46578\,
            I => \N__46566\
        );

    \I__10701\ : Span4Mux_v
    port map (
            O => \N__46575\,
            I => \N__46566\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__46572\,
            I => \N__46563\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46560\
        );

    \I__10698\ : Span4Mux_h
    port map (
            O => \N__46566\,
            I => \N__46555\
        );

    \I__10697\ : Span4Mux_v
    port map (
            O => \N__46563\,
            I => \N__46555\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__46560\,
            I => n20663
        );

    \I__10695\ : Odrv4
    port map (
            O => \N__46555\,
            I => n20663
        );

    \I__10694\ : CascadeMux
    port map (
            O => \N__46550\,
            I => \n12467_cascade_\
        );

    \I__10693\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46544\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46540\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46543\,
            I => \N__46537\
        );

    \I__10690\ : Span4Mux_h
    port map (
            O => \N__46540\,
            I => \N__46532\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__46537\,
            I => \N__46532\
        );

    \I__10688\ : Span4Mux_h
    port map (
            O => \N__46532\,
            I => \N__46529\
        );

    \I__10687\ : Span4Mux_h
    port map (
            O => \N__46529\,
            I => \N__46526\
        );

    \I__10686\ : Odrv4
    port map (
            O => \N__46526\,
            I => n14_adj_1533
        );

    \I__10685\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46518\
        );

    \I__10684\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46515\
        );

    \I__10683\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46512\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46518\,
            I => \N__46509\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46506\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__46512\,
            I => \N__46499\
        );

    \I__10679\ : Span4Mux_v
    port map (
            O => \N__46509\,
            I => \N__46499\
        );

    \I__10678\ : Span4Mux_v
    port map (
            O => \N__46506\,
            I => \N__46499\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__46499\,
            I => data_cntvec_6
        );

    \I__10676\ : InMux
    port map (
            O => \N__46496\,
            I => \N__46493\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__46493\,
            I => \N__46488\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46492\,
            I => \N__46485\
        );

    \I__10673\ : InMux
    port map (
            O => \N__46491\,
            I => \N__46482\
        );

    \I__10672\ : Span4Mux_h
    port map (
            O => \N__46488\,
            I => \N__46479\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__46485\,
            I => \N__46476\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__46482\,
            I => data_cntvec_0
        );

    \I__10669\ : Odrv4
    port map (
            O => \N__46479\,
            I => data_cntvec_0
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__46476\,
            I => data_cntvec_0
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__46469\,
            I => \N__46466\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46462\
        );

    \I__10665\ : CascadeMux
    port map (
            O => \N__46465\,
            I => \N__46458\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__46462\,
            I => \N__46455\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46450\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46450\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__46455\,
            I => req_data_cnt_0
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46450\,
            I => req_data_cnt_0
        );

    \I__10659\ : InMux
    port map (
            O => \N__46445\,
            I => \N__46442\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__46442\,
            I => \N__46439\
        );

    \I__10657\ : Odrv4
    port map (
            O => \N__46439\,
            I => n17
        );

    \I__10656\ : InMux
    port map (
            O => \N__46436\,
            I => \N__46433\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46433\,
            I => \N__46430\
        );

    \I__10654\ : Span4Mux_h
    port map (
            O => \N__46430\,
            I => \N__46427\
        );

    \I__10653\ : Span4Mux_h
    port map (
            O => \N__46427\,
            I => \N__46424\
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__46424\,
            I => n16_adj_1515
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__46421\,
            I => \N__46417\
        );

    \I__10650\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46414\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46411\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46407\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46411\,
            I => \N__46402\
        );

    \I__10646\ : CascadeMux
    port map (
            O => \N__46410\,
            I => \N__46399\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46407\,
            I => \N__46396\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46406\,
            I => \N__46393\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46405\,
            I => \N__46390\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__46402\,
            I => \N__46387\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46399\,
            I => \N__46384\
        );

    \I__10640\ : Span4Mux_v
    port map (
            O => \N__46396\,
            I => \N__46379\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46393\,
            I => \N__46379\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46376\
        );

    \I__10637\ : Span4Mux_h
    port map (
            O => \N__46387\,
            I => \N__46371\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__46384\,
            I => \N__46371\
        );

    \I__10635\ : Span4Mux_v
    port map (
            O => \N__46379\,
            I => \N__46368\
        );

    \I__10634\ : Span4Mux_v
    port map (
            O => \N__46376\,
            I => \N__46362\
        );

    \I__10633\ : Span4Mux_v
    port map (
            O => \N__46371\,
            I => \N__46362\
        );

    \I__10632\ : Span4Mux_h
    port map (
            O => \N__46368\,
            I => \N__46359\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46367\,
            I => \N__46356\
        );

    \I__10630\ : Span4Mux_h
    port map (
            O => \N__46362\,
            I => \N__46352\
        );

    \I__10629\ : Span4Mux_h
    port map (
            O => \N__46359\,
            I => \N__46347\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46347\
        );

    \I__10627\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46344\
        );

    \I__10626\ : Span4Mux_v
    port map (
            O => \N__46352\,
            I => \N__46341\
        );

    \I__10625\ : Span4Mux_v
    port map (
            O => \N__46347\,
            I => \N__46336\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__46344\,
            I => \N__46336\
        );

    \I__10623\ : Odrv4
    port map (
            O => \N__46341\,
            I => comm_buf_0_5
        );

    \I__10622\ : Odrv4
    port map (
            O => \N__46336\,
            I => comm_buf_0_5
        );

    \I__10621\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46328\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__46328\,
            I => \N__46325\
        );

    \I__10619\ : Span4Mux_h
    port map (
            O => \N__46325\,
            I => \N__46320\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46324\,
            I => \N__46315\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46323\,
            I => \N__46315\
        );

    \I__10616\ : Odrv4
    port map (
            O => \N__46320\,
            I => req_data_cnt_6
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__46315\,
            I => req_data_cnt_6
        );

    \I__10614\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46305\
        );

    \I__10613\ : InMux
    port map (
            O => \N__46309\,
            I => \N__46302\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46299\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__46305\,
            I => req_data_cnt_2
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__46302\,
            I => req_data_cnt_2
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__46299\,
            I => req_data_cnt_2
        );

    \I__10608\ : CascadeMux
    port map (
            O => \N__46292\,
            I => \n22208_cascade_\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46289\,
            I => \N__46285\
        );

    \I__10606\ : CascadeMux
    port map (
            O => \N__46288\,
            I => \N__46282\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46285\,
            I => \N__46279\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46282\,
            I => \N__46275\
        );

    \I__10603\ : Span4Mux_v
    port map (
            O => \N__46279\,
            I => \N__46272\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46269\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46275\,
            I => \acadc_skipCount_2\
        );

    \I__10600\ : Odrv4
    port map (
            O => \N__46272\,
            I => \acadc_skipCount_2\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__46269\,
            I => \acadc_skipCount_2\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46262\,
            I => \N__46259\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__46259\,
            I => \N__46256\
        );

    \I__10596\ : Odrv4
    port map (
            O => \N__46256\,
            I => n21959
        );

    \I__10595\ : InMux
    port map (
            O => \N__46253\,
            I => \N__46250\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__46250\,
            I => \N__46247\
        );

    \I__10593\ : Span4Mux_v
    port map (
            O => \N__46247\,
            I => \N__46244\
        );

    \I__10592\ : Odrv4
    port map (
            O => \N__46244\,
            I => comm_buf_3_7
        );

    \I__10591\ : InMux
    port map (
            O => \N__46241\,
            I => \N__46238\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__46238\,
            I => \N__46235\
        );

    \I__10589\ : Span4Mux_v
    port map (
            O => \N__46235\,
            I => \N__46232\
        );

    \I__10588\ : Span4Mux_h
    port map (
            O => \N__46232\,
            I => \N__46229\
        );

    \I__10587\ : Odrv4
    port map (
            O => \N__46229\,
            I => comm_buf_2_7
        );

    \I__10586\ : CascadeMux
    port map (
            O => \N__46226\,
            I => \n2_adj_1581_cascade_\
        );

    \I__10585\ : CEMux
    port map (
            O => \N__46223\,
            I => \N__46220\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46220\,
            I => \N__46215\
        );

    \I__10583\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46209\
        );

    \I__10582\ : CEMux
    port map (
            O => \N__46218\,
            I => \N__46206\
        );

    \I__10581\ : Span4Mux_v
    port map (
            O => \N__46215\,
            I => \N__46202\
        );

    \I__10580\ : CEMux
    port map (
            O => \N__46214\,
            I => \N__46199\
        );

    \I__10579\ : CEMux
    port map (
            O => \N__46213\,
            I => \N__46195\
        );

    \I__10578\ : CEMux
    port map (
            O => \N__46212\,
            I => \N__46192\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__46209\,
            I => \N__46189\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46206\,
            I => \N__46186\
        );

    \I__10575\ : CEMux
    port map (
            O => \N__46205\,
            I => \N__46183\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__46202\,
            I => \N__46178\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__46199\,
            I => \N__46178\
        );

    \I__10572\ : CEMux
    port map (
            O => \N__46198\,
            I => \N__46175\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46195\,
            I => \N__46172\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__46192\,
            I => \N__46169\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__46189\,
            I => \N__46166\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__46186\,
            I => \N__46161\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__46183\,
            I => \N__46161\
        );

    \I__10566\ : Span4Mux_v
    port map (
            O => \N__46178\,
            I => \N__46156\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__46175\,
            I => \N__46156\
        );

    \I__10564\ : Span4Mux_v
    port map (
            O => \N__46172\,
            I => \N__46149\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__46169\,
            I => \N__46149\
        );

    \I__10562\ : Span4Mux_v
    port map (
            O => \N__46166\,
            I => \N__46149\
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__46161\,
            I => n11503
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__46156\,
            I => n11503
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__46149\,
            I => n11503
        );

    \I__10558\ : SRMux
    port map (
            O => \N__46142\,
            I => \N__46137\
        );

    \I__10557\ : SRMux
    port map (
            O => \N__46141\,
            I => \N__46134\
        );

    \I__10556\ : SRMux
    port map (
            O => \N__46140\,
            I => \N__46129\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46137\,
            I => \N__46126\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46123\
        );

    \I__10553\ : SRMux
    port map (
            O => \N__46133\,
            I => \N__46120\
        );

    \I__10552\ : SRMux
    port map (
            O => \N__46132\,
            I => \N__46117\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46112\
        );

    \I__10550\ : Span4Mux_v
    port map (
            O => \N__46126\,
            I => \N__46103\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__46123\,
            I => \N__46103\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__46120\,
            I => \N__46103\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__46117\,
            I => \N__46103\
        );

    \I__10546\ : SRMux
    port map (
            O => \N__46116\,
            I => \N__46100\
        );

    \I__10545\ : SRMux
    port map (
            O => \N__46115\,
            I => \N__46097\
        );

    \I__10544\ : Span4Mux_v
    port map (
            O => \N__46112\,
            I => \N__46094\
        );

    \I__10543\ : Span4Mux_v
    port map (
            O => \N__46103\,
            I => \N__46091\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__46100\,
            I => \N__46088\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__46097\,
            I => \N__46085\
        );

    \I__10540\ : Span4Mux_h
    port map (
            O => \N__46094\,
            I => \N__46080\
        );

    \I__10539\ : Span4Mux_h
    port map (
            O => \N__46091\,
            I => \N__46080\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__46088\,
            I => \N__46077\
        );

    \I__10537\ : Span4Mux_v
    port map (
            O => \N__46085\,
            I => \N__46074\
        );

    \I__10536\ : Odrv4
    port map (
            O => \N__46080\,
            I => n14815
        );

    \I__10535\ : Odrv4
    port map (
            O => \N__46077\,
            I => n14815
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__46074\,
            I => n14815
        );

    \I__10533\ : CascadeMux
    port map (
            O => \N__46067\,
            I => \N__46063\
        );

    \I__10532\ : CascadeMux
    port map (
            O => \N__46066\,
            I => \N__46060\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46063\,
            I => \N__46055\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46052\
        );

    \I__10529\ : InMux
    port map (
            O => \N__46059\,
            I => \N__46049\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__46058\,
            I => \N__46045\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__46055\,
            I => \N__46042\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__46052\,
            I => \N__46038\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__46049\,
            I => \N__46035\
        );

    \I__10524\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46032\
        );

    \I__10523\ : InMux
    port map (
            O => \N__46045\,
            I => \N__46029\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__46042\,
            I => \N__46025\
        );

    \I__10521\ : InMux
    port map (
            O => \N__46041\,
            I => \N__46022\
        );

    \I__10520\ : Span4Mux_h
    port map (
            O => \N__46038\,
            I => \N__46017\
        );

    \I__10519\ : Span4Mux_h
    port map (
            O => \N__46035\,
            I => \N__46017\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__46014\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__46029\,
            I => \N__46011\
        );

    \I__10516\ : CascadeMux
    port map (
            O => \N__46028\,
            I => \N__46008\
        );

    \I__10515\ : Span4Mux_h
    port map (
            O => \N__46025\,
            I => \N__46005\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__46022\,
            I => \N__46002\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__46017\,
            I => \N__45997\
        );

    \I__10512\ : Span4Mux_v
    port map (
            O => \N__46014\,
            I => \N__45997\
        );

    \I__10511\ : Span4Mux_v
    port map (
            O => \N__46011\,
            I => \N__45994\
        );

    \I__10510\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45991\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__46005\,
            I => \N__45986\
        );

    \I__10508\ : Span4Mux_h
    port map (
            O => \N__46002\,
            I => \N__45986\
        );

    \I__10507\ : Sp12to4
    port map (
            O => \N__45997\,
            I => \N__45983\
        );

    \I__10506\ : Sp12to4
    port map (
            O => \N__45994\,
            I => \N__45978\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45991\,
            I => \N__45978\
        );

    \I__10504\ : Span4Mux_v
    port map (
            O => \N__45986\,
            I => \N__45975\
        );

    \I__10503\ : Span12Mux_h
    port map (
            O => \N__45983\,
            I => \N__45970\
        );

    \I__10502\ : Span12Mux_h
    port map (
            O => \N__45978\,
            I => \N__45970\
        );

    \I__10501\ : Odrv4
    port map (
            O => \N__45975\,
            I => comm_buf_0_7
        );

    \I__10500\ : Odrv12
    port map (
            O => \N__45970\,
            I => comm_buf_0_7
        );

    \I__10499\ : InMux
    port map (
            O => \N__45965\,
            I => \N__45962\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__45962\,
            I => n1_adj_1580
        );

    \I__10497\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45956\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45956\,
            I => \N__45953\
        );

    \I__10495\ : Span4Mux_v
    port map (
            O => \N__45953\,
            I => \N__45950\
        );

    \I__10494\ : Span4Mux_h
    port map (
            O => \N__45950\,
            I => \N__45947\
        );

    \I__10493\ : Odrv4
    port map (
            O => \N__45947\,
            I => comm_buf_5_7
        );

    \I__10492\ : InMux
    port map (
            O => \N__45944\,
            I => \N__45941\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__45941\,
            I => \N__45938\
        );

    \I__10490\ : Span4Mux_h
    port map (
            O => \N__45938\,
            I => \N__45935\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__45935\,
            I => comm_buf_4_7
        );

    \I__10488\ : InMux
    port map (
            O => \N__45932\,
            I => \N__45929\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45929\,
            I => n20966
        );

    \I__10486\ : CascadeMux
    port map (
            O => \N__45926\,
            I => \n4_adj_1582_cascade_\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45920\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__45920\,
            I => n21968
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45917\,
            I => \N__45913\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45908\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45913\,
            I => \N__45905\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45902\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45899\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45908\,
            I => \N__45896\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45905\,
            I => \N__45893\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45902\,
            I => \N__45890\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__45899\,
            I => \N__45887\
        );

    \I__10474\ : Span4Mux_v
    port map (
            O => \N__45896\,
            I => \N__45883\
        );

    \I__10473\ : Span4Mux_v
    port map (
            O => \N__45893\,
            I => \N__45880\
        );

    \I__10472\ : Span4Mux_v
    port map (
            O => \N__45890\,
            I => \N__45877\
        );

    \I__10471\ : Span4Mux_h
    port map (
            O => \N__45887\,
            I => \N__45874\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45871\
        );

    \I__10469\ : Sp12to4
    port map (
            O => \N__45883\,
            I => \N__45868\
        );

    \I__10468\ : Span4Mux_v
    port map (
            O => \N__45880\,
            I => \N__45863\
        );

    \I__10467\ : Span4Mux_v
    port map (
            O => \N__45877\,
            I => \N__45863\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__45874\,
            I => comm_buf_1_5
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__45871\,
            I => comm_buf_1_5
        );

    \I__10464\ : Odrv12
    port map (
            O => \N__45868\,
            I => comm_buf_1_5
        );

    \I__10463\ : Odrv4
    port map (
            O => \N__45863\,
            I => comm_buf_1_5
        );

    \I__10462\ : InMux
    port map (
            O => \N__45854\,
            I => \N__45851\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__45851\,
            I => \N__45848\
        );

    \I__10460\ : Span4Mux_h
    port map (
            O => \N__45848\,
            I => \N__45845\
        );

    \I__10459\ : Span4Mux_v
    port map (
            O => \N__45845\,
            I => \N__45842\
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__45842\,
            I => buf_data_iac_9
        );

    \I__10457\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45836\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45836\,
            I => \N__45833\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45833\,
            I => n21270
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__45830\,
            I => \n22241_cascade_\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45827\,
            I => \N__45824\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__45824\,
            I => n8_adj_1576
        );

    \I__10451\ : InMux
    port map (
            O => \N__45821\,
            I => \N__45815\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45820\,
            I => \N__45815\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45815\,
            I => n1272
        );

    \I__10448\ : InMux
    port map (
            O => \N__45812\,
            I => \N__45809\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__45809\,
            I => n20697
        );

    \I__10446\ : InMux
    port map (
            O => \N__45806\,
            I => \N__45803\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45803\,
            I => n4_adj_1614
        );

    \I__10444\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45794\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45794\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45794\,
            I => \N__45791\
        );

    \I__10441\ : Odrv12
    port map (
            O => \N__45791\,
            I => n20668
        );

    \I__10440\ : CEMux
    port map (
            O => \N__45788\,
            I => \N__45785\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45785\,
            I => \N__45782\
        );

    \I__10438\ : Span4Mux_h
    port map (
            O => \N__45782\,
            I => \N__45779\
        );

    \I__10437\ : Span4Mux_v
    port map (
            O => \N__45779\,
            I => \N__45776\
        );

    \I__10436\ : Span4Mux_h
    port map (
            O => \N__45776\,
            I => \N__45773\
        );

    \I__10435\ : Odrv4
    port map (
            O => \N__45773\,
            I => n11866
        );

    \I__10434\ : SRMux
    port map (
            O => \N__45770\,
            I => \N__45767\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45767\,
            I => n14753
        );

    \I__10432\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45761\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__45761\,
            I => \N__45758\
        );

    \I__10430\ : Span4Mux_h
    port map (
            O => \N__45758\,
            I => \N__45755\
        );

    \I__10429\ : Odrv4
    port map (
            O => \N__45755\,
            I => n8_adj_1530
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__45752\,
            I => \n4_adj_1598_cascade_\
        );

    \I__10427\ : CEMux
    port map (
            O => \N__45749\,
            I => \N__45746\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45746\,
            I => n20573
        );

    \I__10425\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45739\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45742\,
            I => \N__45736\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45739\,
            I => \N__45733\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__45736\,
            I => \N__45730\
        );

    \I__10421\ : Span4Mux_h
    port map (
            O => \N__45733\,
            I => \N__45727\
        );

    \I__10420\ : Span12Mux_h
    port map (
            O => \N__45730\,
            I => \N__45724\
        );

    \I__10419\ : Odrv4
    port map (
            O => \N__45727\,
            I => \comm_state_3_N_420_3\
        );

    \I__10418\ : Odrv12
    port map (
            O => \N__45724\,
            I => \comm_state_3_N_420_3\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__45719\,
            I => \n1272_cascade_\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45713\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__45713\,
            I => \N__45710\
        );

    \I__10414\ : Span4Mux_v
    port map (
            O => \N__45710\,
            I => \N__45707\
        );

    \I__10413\ : Odrv4
    port map (
            O => \N__45707\,
            I => comm_buf_4_5
        );

    \I__10412\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45701\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45701\,
            I => n22175
        );

    \I__10410\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45695\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__45695\,
            I => n20551
        );

    \I__10408\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45689\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__45689\,
            I => \N__45686\
        );

    \I__10406\ : Odrv4
    port map (
            O => \N__45686\,
            I => n11420
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__45683\,
            I => \n20551_cascade_\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45677\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__10402\ : Odrv4
    port map (
            O => \N__45674\,
            I => n20717
        );

    \I__10401\ : CEMux
    port map (
            O => \N__45671\,
            I => \N__45668\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10399\ : Span4Mux_h
    port map (
            O => \N__45665\,
            I => \N__45662\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__45662\,
            I => n20575
        );

    \I__10397\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45656\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__45656\,
            I => \N__45653\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__45653\,
            I => \N__45650\
        );

    \I__10394\ : Span4Mux_h
    port map (
            O => \N__45650\,
            I => \N__45647\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__45647\,
            I => n20962
        );

    \I__10392\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45640\
        );

    \I__10391\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45637\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45633\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45637\,
            I => \N__45630\
        );

    \I__10388\ : CascadeMux
    port map (
            O => \N__45636\,
            I => \N__45627\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__45633\,
            I => \N__45622\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__45630\,
            I => \N__45622\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45619\
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__45622\,
            I => n14545
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__45619\,
            I => n14545
        );

    \I__10382\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45611\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__45611\,
            I => n22238
        );

    \I__10380\ : CascadeMux
    port map (
            O => \N__45608\,
            I => \n2_adj_1575_cascade_\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45602\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45602\,
            I => \N__45599\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__10376\ : Odrv4
    port map (
            O => \N__45596\,
            I => comm_buf_2_1
        );

    \I__10375\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45590\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__45590\,
            I => \N__45587\
        );

    \I__10373\ : Span4Mux_h
    port map (
            O => \N__45587\,
            I => \N__45584\
        );

    \I__10372\ : Odrv4
    port map (
            O => \N__45584\,
            I => comm_buf_3_1
        );

    \I__10371\ : CascadeMux
    port map (
            O => \N__45581\,
            I => \N__45578\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45573\
        );

    \I__10369\ : CascadeMux
    port map (
            O => \N__45577\,
            I => \N__45570\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__45576\,
            I => \N__45567\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__45573\,
            I => \N__45563\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45560\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45557\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45553\
        );

    \I__10363\ : Span4Mux_v
    port map (
            O => \N__45563\,
            I => \N__45546\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__45560\,
            I => \N__45546\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__45557\,
            I => \N__45546\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45541\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45538\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__45546\,
            I => \N__45533\
        );

    \I__10357\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45530\
        );

    \I__10356\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45527\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__45541\,
            I => \N__45522\
        );

    \I__10354\ : Span4Mux_v
    port map (
            O => \N__45538\,
            I => \N__45522\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45518\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45515\
        );

    \I__10351\ : Span4Mux_v
    port map (
            O => \N__45533\,
            I => \N__45510\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45530\,
            I => \N__45510\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45527\,
            I => \N__45505\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__45522\,
            I => \N__45505\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45521\,
            I => \N__45502\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__45518\,
            I => \N__45499\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__45515\,
            I => \N__45496\
        );

    \I__10344\ : Span4Mux_v
    port map (
            O => \N__45510\,
            I => \N__45493\
        );

    \I__10343\ : Sp12to4
    port map (
            O => \N__45505\,
            I => \N__45488\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__45502\,
            I => \N__45488\
        );

    \I__10341\ : Span4Mux_h
    port map (
            O => \N__45499\,
            I => \N__45485\
        );

    \I__10340\ : Span12Mux_v
    port map (
            O => \N__45496\,
            I => \N__45482\
        );

    \I__10339\ : Sp12to4
    port map (
            O => \N__45493\,
            I => \N__45477\
        );

    \I__10338\ : Span12Mux_v
    port map (
            O => \N__45488\,
            I => \N__45477\
        );

    \I__10337\ : Odrv4
    port map (
            O => \N__45485\,
            I => comm_buf_0_1
        );

    \I__10336\ : Odrv12
    port map (
            O => \N__45482\,
            I => comm_buf_0_1
        );

    \I__10335\ : Odrv12
    port map (
            O => \N__45477\,
            I => comm_buf_0_1
        );

    \I__10334\ : CascadeMux
    port map (
            O => \N__45470\,
            I => \n22052_cascade_\
        );

    \I__10333\ : CascadeMux
    port map (
            O => \N__45467\,
            I => \N__45464\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45464\,
            I => \N__45461\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45461\,
            I => \N__45458\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__45458\,
            I => \N__45450\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45441\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45441\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45441\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45441\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45438\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__45450\,
            I => \N__45435\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__45441\,
            I => \N__45432\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45438\,
            I => \N__45429\
        );

    \I__10321\ : Span4Mux_h
    port map (
            O => \N__45435\,
            I => \N__45424\
        );

    \I__10320\ : Span4Mux_h
    port map (
            O => \N__45432\,
            I => \N__45424\
        );

    \I__10319\ : Span4Mux_v
    port map (
            O => \N__45429\,
            I => \N__45421\
        );

    \I__10318\ : Span4Mux_v
    port map (
            O => \N__45424\,
            I => \N__45418\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__45421\,
            I => comm_buf_1_1
        );

    \I__10316\ : Odrv4
    port map (
            O => \N__45418\,
            I => comm_buf_1_1
        );

    \I__10315\ : InMux
    port map (
            O => \N__45413\,
            I => \N__45410\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__45410\,
            I => n20807
        );

    \I__10313\ : CascadeMux
    port map (
            O => \N__45407\,
            I => \n22055_cascade_\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45401\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45401\,
            I => \N__45398\
        );

    \I__10310\ : Span4Mux_h
    port map (
            O => \N__45398\,
            I => \N__45395\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__45395\,
            I => comm_buf_5_5
        );

    \I__10308\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45389\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__45389\,
            I => \N__45386\
        );

    \I__10306\ : Odrv12
    port map (
            O => \N__45386\,
            I => comm_buf_3_5
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__45383\,
            I => \n17404_cascade_\
        );

    \I__10304\ : CascadeMux
    port map (
            O => \N__45380\,
            I => \n20951_cascade_\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45373\
        );

    \I__10302\ : CascadeMux
    port map (
            O => \N__45376\,
            I => \N__45369\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__45373\,
            I => \N__45366\
        );

    \I__10300\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45359\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45369\,
            I => \N__45356\
        );

    \I__10298\ : Span4Mux_v
    port map (
            O => \N__45366\,
            I => \N__45353\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45365\,
            I => \N__45350\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45347\
        );

    \I__10295\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45344\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45341\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__45359\,
            I => \N__45338\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__45356\,
            I => \N__45335\
        );

    \I__10291\ : Span4Mux_v
    port map (
            O => \N__45353\,
            I => \N__45330\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__45350\,
            I => \N__45330\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45347\,
            I => \N__45323\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45344\,
            I => \N__45323\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45323\
        );

    \I__10286\ : Span4Mux_v
    port map (
            O => \N__45338\,
            I => \N__45318\
        );

    \I__10285\ : Span4Mux_v
    port map (
            O => \N__45335\,
            I => \N__45315\
        );

    \I__10284\ : Span4Mux_h
    port map (
            O => \N__45330\,
            I => \N__45312\
        );

    \I__10283\ : Span4Mux_v
    port map (
            O => \N__45323\,
            I => \N__45309\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45306\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45303\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__45318\,
            I => comm_rx_buf_1
        );

    \I__10279\ : Odrv4
    port map (
            O => \N__45315\,
            I => comm_rx_buf_1
        );

    \I__10278\ : Odrv4
    port map (
            O => \N__45312\,
            I => comm_rx_buf_1
        );

    \I__10277\ : Odrv4
    port map (
            O => \N__45309\,
            I => comm_rx_buf_1
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__45306\,
            I => comm_rx_buf_1
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__45303\,
            I => comm_rx_buf_1
        );

    \I__10274\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45286\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45289\,
            I => \N__45283\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__45286\,
            I => comm_buf_6_1
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__45283\,
            I => comm_buf_6_1
        );

    \I__10270\ : IoInMux
    port map (
            O => \N__45278\,
            I => \N__45275\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__45275\,
            I => \N__45272\
        );

    \I__10268\ : Span4Mux_s3_v
    port map (
            O => \N__45272\,
            I => \N__45269\
        );

    \I__10267\ : Span4Mux_v
    port map (
            O => \N__45269\,
            I => \N__45266\
        );

    \I__10266\ : Sp12to4
    port map (
            O => \N__45266\,
            I => \N__45263\
        );

    \I__10265\ : Odrv12
    port map (
            O => \N__45263\,
            I => \DDS_CS\
        );

    \I__10264\ : CEMux
    port map (
            O => \N__45260\,
            I => \N__45257\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__45257\,
            I => \N__45254\
        );

    \I__10262\ : Span4Mux_v
    port map (
            O => \N__45254\,
            I => \N__45251\
        );

    \I__10261\ : Span4Mux_h
    port map (
            O => \N__45251\,
            I => \N__45248\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__45248\,
            I => \SIG_DDS.n9_adj_1394\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45242\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45242\,
            I => \N__45239\
        );

    \I__10257\ : Span4Mux_h
    port map (
            O => \N__45239\,
            I => \N__45236\
        );

    \I__10256\ : Odrv4
    port map (
            O => \N__45236\,
            I => buf_data_iac_20
        );

    \I__10255\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45230\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__45230\,
            I => \N__45227\
        );

    \I__10253\ : Span4Mux_h
    port map (
            O => \N__45227\,
            I => \N__45224\
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__45224\,
            I => n20984
        );

    \I__10251\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45218\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__45218\,
            I => n17738
        );

    \I__10249\ : CascadeMux
    port map (
            O => \N__45215\,
            I => \N__45212\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45209\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__45209\,
            I => n14146
        );

    \I__10246\ : CascadeMux
    port map (
            O => \N__45206\,
            I => \N__45202\
        );

    \I__10245\ : CascadeMux
    port map (
            O => \N__45205\,
            I => \N__45198\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45195\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45188\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45198\,
            I => \N__45188\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__45195\,
            I => \N__45184\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45181\
        );

    \I__10239\ : InMux
    port map (
            O => \N__45193\,
            I => \N__45178\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__45188\,
            I => \N__45175\
        );

    \I__10237\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45172\
        );

    \I__10236\ : Span4Mux_v
    port map (
            O => \N__45184\,
            I => \N__45167\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45167\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__45178\,
            I => \N__45162\
        );

    \I__10233\ : Span4Mux_h
    port map (
            O => \N__45175\,
            I => \N__45162\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__45172\,
            I => \N__45159\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__45167\,
            I => \N__45156\
        );

    \I__10230\ : Span4Mux_v
    port map (
            O => \N__45162\,
            I => \N__45153\
        );

    \I__10229\ : Span4Mux_h
    port map (
            O => \N__45159\,
            I => \N__45150\
        );

    \I__10228\ : Sp12to4
    port map (
            O => \N__45156\,
            I => \N__45147\
        );

    \I__10227\ : Span4Mux_h
    port map (
            O => \N__45153\,
            I => \N__45144\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__45150\,
            I => \comm_state_3_N_436_2\
        );

    \I__10225\ : Odrv12
    port map (
            O => \N__45147\,
            I => \comm_state_3_N_436_2\
        );

    \I__10224\ : Odrv4
    port map (
            O => \N__45144\,
            I => \comm_state_3_N_436_2\
        );

    \I__10223\ : CascadeMux
    port map (
            O => \N__45137\,
            I => \n15_cascade_\
        );

    \I__10222\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45131\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__45131\,
            I => n12_adj_1649
        );

    \I__10220\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45125\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__45125\,
            I => \N__45122\
        );

    \I__10218\ : Span4Mux_h
    port map (
            O => \N__45122\,
            I => \N__45119\
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__45119\,
            I => comm_buf_4_1
        );

    \I__10216\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45113\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45110\
        );

    \I__10214\ : Span4Mux_v
    port map (
            O => \N__45110\,
            I => \N__45107\
        );

    \I__10213\ : Span4Mux_h
    port map (
            O => \N__45107\,
            I => \N__45104\
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__45104\,
            I => comm_buf_5_1
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__45101\,
            I => \n4_adj_1595_cascade_\
        );

    \I__10210\ : InMux
    port map (
            O => \N__45098\,
            I => \N__45094\
        );

    \I__10209\ : InMux
    port map (
            O => \N__45097\,
            I => \N__45091\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__45094\,
            I => \N__45087\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__45091\,
            I => \N__45075\
        );

    \I__10206\ : ClkMux
    port map (
            O => \N__45090\,
            I => \N__45035\
        );

    \I__10205\ : Glb2LocalMux
    port map (
            O => \N__45087\,
            I => \N__45035\
        );

    \I__10204\ : ClkMux
    port map (
            O => \N__45086\,
            I => \N__45035\
        );

    \I__10203\ : ClkMux
    port map (
            O => \N__45085\,
            I => \N__45035\
        );

    \I__10202\ : ClkMux
    port map (
            O => \N__45084\,
            I => \N__45035\
        );

    \I__10201\ : ClkMux
    port map (
            O => \N__45083\,
            I => \N__45035\
        );

    \I__10200\ : ClkMux
    port map (
            O => \N__45082\,
            I => \N__45035\
        );

    \I__10199\ : ClkMux
    port map (
            O => \N__45081\,
            I => \N__45035\
        );

    \I__10198\ : ClkMux
    port map (
            O => \N__45080\,
            I => \N__45035\
        );

    \I__10197\ : ClkMux
    port map (
            O => \N__45079\,
            I => \N__45035\
        );

    \I__10196\ : ClkMux
    port map (
            O => \N__45078\,
            I => \N__45035\
        );

    \I__10195\ : Glb2LocalMux
    port map (
            O => \N__45075\,
            I => \N__45035\
        );

    \I__10194\ : ClkMux
    port map (
            O => \N__45074\,
            I => \N__45035\
        );

    \I__10193\ : ClkMux
    port map (
            O => \N__45073\,
            I => \N__45035\
        );

    \I__10192\ : ClkMux
    port map (
            O => \N__45072\,
            I => \N__45035\
        );

    \I__10191\ : ClkMux
    port map (
            O => \N__45071\,
            I => \N__45035\
        );

    \I__10190\ : ClkMux
    port map (
            O => \N__45070\,
            I => \N__45035\
        );

    \I__10189\ : GlobalMux
    port map (
            O => \N__45035\,
            I => \clk_16MHz\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45032\,
            I => \N__45029\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__45029\,
            I => \N__45025\
        );

    \I__10186\ : InMux
    port map (
            O => \N__45028\,
            I => \N__45022\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__45025\,
            I => dds0_mclk
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__45022\,
            I => dds0_mclk
        );

    \I__10183\ : InMux
    port map (
            O => \N__45017\,
            I => \N__45013\
        );

    \I__10182\ : InMux
    port map (
            O => \N__45016\,
            I => \N__45009\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__45013\,
            I => \N__45006\
        );

    \I__10180\ : CascadeMux
    port map (
            O => \N__45012\,
            I => \N__45003\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__45000\
        );

    \I__10178\ : Span4Mux_h
    port map (
            O => \N__45006\,
            I => \N__44997\
        );

    \I__10177\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44994\
        );

    \I__10176\ : Span12Mux_h
    port map (
            O => \N__45000\,
            I => \N__44989\
        );

    \I__10175\ : Sp12to4
    port map (
            O => \N__44997\,
            I => \N__44989\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44994\,
            I => buf_control_6
        );

    \I__10173\ : Odrv12
    port map (
            O => \N__44989\,
            I => buf_control_6
        );

    \I__10172\ : IoInMux
    port map (
            O => \N__44984\,
            I => \N__44981\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44981\,
            I => \N__44978\
        );

    \I__10170\ : Span4Mux_s0_v
    port map (
            O => \N__44978\,
            I => \N__44975\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__44975\,
            I => \N__44972\
        );

    \I__10168\ : Sp12to4
    port map (
            O => \N__44972\,
            I => \N__44969\
        );

    \I__10167\ : Span12Mux_h
    port map (
            O => \N__44969\,
            I => \N__44966\
        );

    \I__10166\ : Odrv12
    port map (
            O => \N__44966\,
            I => \DDS_MCLK\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44963\,
            I => \N__44960\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44960\,
            I => \N__44956\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44953\
        );

    \I__10162\ : Span4Mux_h
    port map (
            O => \N__44956\,
            I => \N__44950\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44946\
        );

    \I__10160\ : Span4Mux_h
    port map (
            O => \N__44950\,
            I => \N__44943\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44940\
        );

    \I__10158\ : Span12Mux_h
    port map (
            O => \N__44946\,
            I => \N__44937\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__44943\,
            I => \N__44934\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44940\,
            I => buf_adcdata_iac_15
        );

    \I__10155\ : Odrv12
    port map (
            O => \N__44937\,
            I => buf_adcdata_iac_15
        );

    \I__10154\ : Odrv4
    port map (
            O => \N__44934\,
            I => buf_adcdata_iac_15
        );

    \I__10153\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44924\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__44924\,
            I => n16_adj_1503
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__44921\,
            I => \N__44918\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44918\,
            I => \N__44915\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__44915\,
            I => \N__44912\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__44912\,
            I => \N__44909\
        );

    \I__10147\ : Odrv4
    port map (
            O => \N__44909\,
            I => n20797
        );

    \I__10146\ : InMux
    port map (
            O => \N__44906\,
            I => \N__44902\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44905\,
            I => \N__44899\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44902\,
            I => \N__44894\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44891\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44886\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44886\
        );

    \I__10140\ : Odrv12
    port map (
            O => \N__44894\,
            I => eis_stop
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__44891\,
            I => eis_stop
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44886\,
            I => eis_stop
        );

    \I__10137\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44876\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44876\,
            I => \N__44873\
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__44873\,
            I => n22034
        );

    \I__10134\ : CascadeMux
    port map (
            O => \N__44870\,
            I => \N__44866\
        );

    \I__10133\ : CascadeMux
    port map (
            O => \N__44869\,
            I => \N__44863\
        );

    \I__10132\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44854\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44854\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44854\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44861\,
            I => \N__44851\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44854\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44851\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__10126\ : CascadeMux
    port map (
            O => \N__44846\,
            I => \N__44841\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44845\,
            I => \N__44836\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44836\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44833\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44836\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44833\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44828\,
            I => \N__44824\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44821\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44824\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44821\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44816\,
            I => \N__44812\
        );

    \I__10115\ : CascadeMux
    port map (
            O => \N__44815\,
            I => \N__44808\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44805\
        );

    \I__10113\ : CascadeMux
    port map (
            O => \N__44811\,
            I => \N__44802\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44808\,
            I => \N__44799\
        );

    \I__10111\ : Span4Mux_v
    port map (
            O => \N__44805\,
            I => \N__44796\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44793\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44799\,
            I => \N__44790\
        );

    \I__10108\ : Span4Mux_h
    port map (
            O => \N__44796\,
            I => \N__44784\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44793\,
            I => \N__44784\
        );

    \I__10106\ : Span4Mux_h
    port map (
            O => \N__44790\,
            I => \N__44781\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44778\
        );

    \I__10104\ : Span4Mux_h
    port map (
            O => \N__44784\,
            I => \N__44775\
        );

    \I__10103\ : Span4Mux_h
    port map (
            O => \N__44781\,
            I => \N__44772\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44778\,
            I => trig_dds0
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__44775\,
            I => trig_dds0
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__44772\,
            I => trig_dds0
        );

    \I__10099\ : SRMux
    port map (
            O => \N__44765\,
            I => \N__44761\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44758\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44761\,
            I => n14900
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44758\,
            I => n14900
        );

    \I__10095\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44742\
        );

    \I__10094\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44742\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44742\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44750\,
            I => \N__44737\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44737\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44742\,
            I => bit_cnt_0
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44737\,
            I => bit_cnt_0
        );

    \I__10088\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44729\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44729\,
            I => \N__44725\
        );

    \I__10086\ : CascadeMux
    port map (
            O => \N__44728\,
            I => \N__44722\
        );

    \I__10085\ : Span4Mux_v
    port map (
            O => \N__44725\,
            I => \N__44719\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44716\
        );

    \I__10083\ : Span4Mux_h
    port map (
            O => \N__44719\,
            I => \N__44713\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__44716\,
            I => \N__44710\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__44713\,
            I => tmp_buf_15
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__44710\,
            I => tmp_buf_15
        );

    \I__10079\ : IoInMux
    port map (
            O => \N__44705\,
            I => \N__44702\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__44702\,
            I => \N__44699\
        );

    \I__10077\ : Span4Mux_s1_v
    port map (
            O => \N__44699\,
            I => \N__44696\
        );

    \I__10076\ : Sp12to4
    port map (
            O => \N__44696\,
            I => \N__44693\
        );

    \I__10075\ : Span12Mux_h
    port map (
            O => \N__44693\,
            I => \N__44689\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44692\,
            I => \N__44686\
        );

    \I__10073\ : Odrv12
    port map (
            O => \N__44689\,
            I => \DDS_MOSI\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__44686\,
            I => \DDS_MOSI\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44681\,
            I => \N__44678\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__44678\,
            I => \N__44675\
        );

    \I__10069\ : Span4Mux_h
    port map (
            O => \N__44675\,
            I => \N__44672\
        );

    \I__10068\ : Span4Mux_h
    port map (
            O => \N__44672\,
            I => \N__44669\
        );

    \I__10067\ : Odrv4
    port map (
            O => \N__44669\,
            I => n22226
        );

    \I__10066\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44663\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__44663\,
            I => n22229
        );

    \I__10064\ : IoInMux
    port map (
            O => \N__44660\,
            I => \N__44657\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__44657\,
            I => \N__44654\
        );

    \I__10062\ : Span4Mux_s0_v
    port map (
            O => \N__44654\,
            I => \N__44650\
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__44653\,
            I => \N__44647\
        );

    \I__10060\ : Span4Mux_v
    port map (
            O => \N__44650\,
            I => \N__44644\
        );

    \I__10059\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44640\
        );

    \I__10058\ : Sp12to4
    port map (
            O => \N__44644\,
            I => \N__44637\
        );

    \I__10057\ : CascadeMux
    port map (
            O => \N__44643\,
            I => \N__44634\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__44640\,
            I => \N__44631\
        );

    \I__10055\ : Span12Mux_h
    port map (
            O => \N__44637\,
            I => \N__44628\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44625\
        );

    \I__10053\ : Span4Mux_h
    port map (
            O => \N__44631\,
            I => \N__44622\
        );

    \I__10052\ : Odrv12
    port map (
            O => \N__44628\,
            I => \DDS_RNG_0\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44625\,
            I => \DDS_RNG_0\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__44622\,
            I => \DDS_RNG_0\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44615\,
            I => \N__44612\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__44612\,
            I => \N__44609\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__44609\,
            I => \N__44604\
        );

    \I__10046\ : InMux
    port map (
            O => \N__44608\,
            I => \N__44599\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44599\
        );

    \I__10044\ : Odrv4
    port map (
            O => \N__44604\,
            I => \acadc_skipCount_9\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__44599\,
            I => \acadc_skipCount_9\
        );

    \I__10042\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44591\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__44591\,
            I => n22037
        );

    \I__10040\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44583\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44587\,
            I => \N__44580\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44577\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__44583\,
            I => \N__44572\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44580\,
            I => \N__44572\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44577\,
            I => buf_dds1_7
        );

    \I__10034\ : Odrv12
    port map (
            O => \N__44572\,
            I => buf_dds1_7
        );

    \I__10033\ : InMux
    port map (
            O => \N__44567\,
            I => \N__44564\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44559\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44556\
        );

    \I__10030\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44553\
        );

    \I__10029\ : Span4Mux_v
    port map (
            O => \N__44559\,
            I => \N__44550\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44556\,
            I => \N__44547\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__44553\,
            I => buf_dds0_7
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__44550\,
            I => buf_dds0_7
        );

    \I__10025\ : Odrv12
    port map (
            O => \N__44547\,
            I => buf_dds0_7
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__44540\,
            I => \N__44537\
        );

    \I__10023\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44533\
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__44536\,
            I => \N__44530\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44533\,
            I => \N__44526\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44523\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44529\,
            I => \N__44520\
        );

    \I__10018\ : Span4Mux_h
    port map (
            O => \N__44526\,
            I => \N__44517\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__44523\,
            I => \N__44514\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__44520\,
            I => req_data_cnt_11
        );

    \I__10015\ : Odrv4
    port map (
            O => \N__44517\,
            I => req_data_cnt_11
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__44514\,
            I => req_data_cnt_11
        );

    \I__10013\ : InMux
    port map (
            O => \N__44507\,
            I => \N__44504\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44504\,
            I => n23_adj_1540
        );

    \I__10011\ : InMux
    port map (
            O => \N__44501\,
            I => \N__44498\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__44498\,
            I => \N__44495\
        );

    \I__10009\ : Sp12to4
    port map (
            O => \N__44495\,
            I => \N__44492\
        );

    \I__10008\ : Odrv12
    port map (
            O => \N__44492\,
            I => n20836
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__44489\,
            I => \N__44485\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44482\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44479\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44482\,
            I => \N__44474\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44479\,
            I => \N__44471\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44468\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44464\
        );

    \I__10000\ : Span4Mux_v
    port map (
            O => \N__44474\,
            I => \N__44457\
        );

    \I__9999\ : Span4Mux_v
    port map (
            O => \N__44471\,
            I => \N__44457\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44468\,
            I => \N__44457\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44467\,
            I => \N__44454\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__44464\,
            I => \N__44451\
        );

    \I__9995\ : Span4Mux_h
    port map (
            O => \N__44457\,
            I => \N__44448\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44454\,
            I => n14_adj_1545
        );

    \I__9993\ : Odrv4
    port map (
            O => \N__44451\,
            I => n14_adj_1545
        );

    \I__9992\ : Odrv4
    port map (
            O => \N__44448\,
            I => n14_adj_1545
        );

    \I__9991\ : InMux
    port map (
            O => \N__44441\,
            I => \N__44435\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__44440\,
            I => \N__44431\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44439\,
            I => \N__44426\
        );

    \I__9988\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44423\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44420\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44415\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44415\
        );

    \I__9984\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44410\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44429\,
            I => \N__44410\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__44426\,
            I => \N__44405\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44405\
        );

    \I__9980\ : Span4Mux_h
    port map (
            O => \N__44420\,
            I => \N__44402\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44399\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44410\,
            I => \N__44396\
        );

    \I__9977\ : Span4Mux_h
    port map (
            O => \N__44405\,
            I => \N__44393\
        );

    \I__9976\ : Span4Mux_h
    port map (
            O => \N__44402\,
            I => \N__44390\
        );

    \I__9975\ : Span4Mux_h
    port map (
            O => \N__44399\,
            I => \N__44387\
        );

    \I__9974\ : Span4Mux_v
    port map (
            O => \N__44396\,
            I => \N__44382\
        );

    \I__9973\ : Span4Mux_v
    port map (
            O => \N__44393\,
            I => \N__44382\
        );

    \I__9972\ : Odrv4
    port map (
            O => \N__44390\,
            I => n11931
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__44387\,
            I => n11931
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__44382\,
            I => n11931
        );

    \I__9969\ : CascadeMux
    port map (
            O => \N__44375\,
            I => \n21073_cascade_\
        );

    \I__9968\ : CascadeMux
    port map (
            O => \N__44372\,
            I => \n21072_cascade_\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44369\,
            I => \N__44366\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__44366\,
            I => n23
        );

    \I__9965\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44360\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__44360\,
            I => n21_adj_1521
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__44357\,
            I => \n22_adj_1568_cascade_\
        );

    \I__9962\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__44351\,
            I => n30_adj_1641
        );

    \I__9960\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44344\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__44347\,
            I => \N__44341\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__44344\,
            I => \N__44338\
        );

    \I__9957\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44335\
        );

    \I__9956\ : Span4Mux_h
    port map (
            O => \N__44338\,
            I => \N__44332\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44335\,
            I => data_idxvec_9
        );

    \I__9954\ : Odrv4
    port map (
            O => \N__44332\,
            I => data_idxvec_9
        );

    \I__9953\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44324\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__44324\,
            I => \N__44321\
        );

    \I__9951\ : Span4Mux_h
    port map (
            O => \N__44321\,
            I => \N__44318\
        );

    \I__9950\ : Span4Mux_h
    port map (
            O => \N__44318\,
            I => \N__44315\
        );

    \I__9949\ : Odrv4
    port map (
            O => \N__44315\,
            I => buf_data_iac_17
        );

    \I__9948\ : CascadeMux
    port map (
            O => \N__44312\,
            I => \n20812_cascade_\
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__44309\,
            I => \N__44304\
        );

    \I__9946\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44298\
        );

    \I__9945\ : InMux
    port map (
            O => \N__44307\,
            I => \N__44295\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44304\,
            I => \N__44292\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__44303\,
            I => \N__44288\
        );

    \I__9942\ : CascadeMux
    port map (
            O => \N__44302\,
            I => \N__44285\
        );

    \I__9941\ : CascadeMux
    port map (
            O => \N__44301\,
            I => \N__44282\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44278\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44295\,
            I => \N__44275\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__44292\,
            I => \N__44272\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44269\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44288\,
            I => \N__44266\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44285\,
            I => \N__44263\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44260\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44281\,
            I => \N__44256\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__44278\,
            I => \N__44253\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__44275\,
            I => \N__44248\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__44272\,
            I => \N__44248\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44269\,
            I => \N__44245\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__44266\,
            I => \N__44242\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__44263\,
            I => \N__44239\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__44260\,
            I => \N__44236\
        );

    \I__9925\ : InMux
    port map (
            O => \N__44259\,
            I => \N__44233\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__44256\,
            I => \N__44228\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__44253\,
            I => \N__44228\
        );

    \I__9922\ : Span4Mux_v
    port map (
            O => \N__44248\,
            I => \N__44223\
        );

    \I__9921\ : Span4Mux_h
    port map (
            O => \N__44245\,
            I => \N__44223\
        );

    \I__9920\ : Span4Mux_v
    port map (
            O => \N__44242\,
            I => \N__44220\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__44239\,
            I => \N__44215\
        );

    \I__9918\ : Span4Mux_v
    port map (
            O => \N__44236\,
            I => \N__44215\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__44233\,
            I => \N__44208\
        );

    \I__9916\ : Span4Mux_h
    port map (
            O => \N__44228\,
            I => \N__44208\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__44223\,
            I => \N__44208\
        );

    \I__9914\ : Odrv4
    port map (
            O => \N__44220\,
            I => comm_buf_0_3
        );

    \I__9913\ : Odrv4
    port map (
            O => \N__44215\,
            I => comm_buf_0_3
        );

    \I__9912\ : Odrv4
    port map (
            O => \N__44208\,
            I => comm_buf_0_3
        );

    \I__9911\ : IoInMux
    port map (
            O => \N__44201\,
            I => \N__44198\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44194\
        );

    \I__9909\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44190\
        );

    \I__9908\ : Span12Mux_s3_v
    port map (
            O => \N__44194\,
            I => \N__44187\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44184\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__44190\,
            I => \N__44181\
        );

    \I__9905\ : Odrv12
    port map (
            O => \N__44187\,
            I => \SELIRNG1\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__44184\,
            I => \SELIRNG1\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__44181\,
            I => \SELIRNG1\
        );

    \I__9902\ : CascadeMux
    port map (
            O => \N__44174\,
            I => \N__44170\
        );

    \I__9901\ : InMux
    port map (
            O => \N__44173\,
            I => \N__44165\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44162\
        );

    \I__9899\ : CascadeMux
    port map (
            O => \N__44169\,
            I => \N__44159\
        );

    \I__9898\ : CascadeMux
    port map (
            O => \N__44168\,
            I => \N__44156\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44165\,
            I => \N__44152\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44149\
        );

    \I__9895\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44146\
        );

    \I__9894\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44143\
        );

    \I__9893\ : InMux
    port map (
            O => \N__44155\,
            I => \N__44140\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__44152\,
            I => \N__44136\
        );

    \I__9891\ : Span4Mux_v
    port map (
            O => \N__44149\,
            I => \N__44133\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__44146\,
            I => \N__44128\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44128\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__44140\,
            I => \N__44124\
        );

    \I__9887\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44121\
        );

    \I__9886\ : Span4Mux_h
    port map (
            O => \N__44136\,
            I => \N__44113\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__44133\,
            I => \N__44113\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__44128\,
            I => \N__44113\
        );

    \I__9883\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44110\
        );

    \I__9882\ : Span4Mux_h
    port map (
            O => \N__44124\,
            I => \N__44105\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__44121\,
            I => \N__44105\
        );

    \I__9880\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44102\
        );

    \I__9879\ : Span4Mux_v
    port map (
            O => \N__44113\,
            I => \N__44099\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__44110\,
            I => \N__44094\
        );

    \I__9877\ : Span4Mux_v
    port map (
            O => \N__44105\,
            I => \N__44094\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44091\
        );

    \I__9875\ : Span4Mux_v
    port map (
            O => \N__44099\,
            I => \N__44088\
        );

    \I__9874\ : Span4Mux_v
    port map (
            O => \N__44094\,
            I => \N__44085\
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__44091\,
            I => comm_buf_0_4
        );

    \I__9872\ : Odrv4
    port map (
            O => \N__44088\,
            I => comm_buf_0_4
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__44085\,
            I => comm_buf_0_4
        );

    \I__9870\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44074\
        );

    \I__9869\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44071\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__44074\,
            I => \N__44068\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__44071\,
            I => \N__44065\
        );

    \I__9866\ : Span4Mux_v
    port map (
            O => \N__44068\,
            I => \N__44062\
        );

    \I__9865\ : Span12Mux_h
    port map (
            O => \N__44065\,
            I => \N__44059\
        );

    \I__9864\ : Odrv4
    port map (
            O => \N__44062\,
            I => n14_adj_1571
        );

    \I__9863\ : Odrv12
    port map (
            O => \N__44059\,
            I => n14_adj_1571
        );

    \I__9862\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44051\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__44051\,
            I => \N__44047\
        );

    \I__9860\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44044\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44041\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__44044\,
            I => \N__44038\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__44041\,
            I => \N__44035\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__44038\,
            I => \N__44032\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__44035\,
            I => \N__44029\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__44032\,
            I => n14_adj_1549
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__44029\,
            I => n14_adj_1549
        );

    \I__9852\ : InMux
    port map (
            O => \N__44024\,
            I => \N__44021\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__44021\,
            I => n20814
        );

    \I__9850\ : InMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__44015\,
            I => \N__44012\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__44009\,
            I => n22025
        );

    \I__9846\ : CascadeMux
    port map (
            O => \N__44006\,
            I => \n22232_cascade_\
        );

    \I__9845\ : InMux
    port map (
            O => \N__44003\,
            I => \N__44000\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__44000\,
            I => \N__43997\
        );

    \I__9843\ : Span12Mux_v
    port map (
            O => \N__43997\,
            I => \N__43994\
        );

    \I__9842\ : Odrv12
    port map (
            O => \N__43994\,
            I => n22235
        );

    \I__9841\ : InMux
    port map (
            O => \N__43991\,
            I => \N__43988\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__43988\,
            I => \N__43985\
        );

    \I__9839\ : Span4Mux_v
    port map (
            O => \N__43985\,
            I => \N__43982\
        );

    \I__9838\ : Sp12to4
    port map (
            O => \N__43982\,
            I => \N__43979\
        );

    \I__9837\ : Span12Mux_h
    port map (
            O => \N__43979\,
            I => \N__43975\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43978\,
            I => \N__43972\
        );

    \I__9835\ : Odrv12
    port map (
            O => \N__43975\,
            I => buf_adcdata_vdc_17
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__43972\,
            I => buf_adcdata_vdc_17
        );

    \I__9833\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43964\,
            I => \N__43961\
        );

    \I__9831\ : Span4Mux_h
    port map (
            O => \N__43961\,
            I => \N__43957\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__43960\,
            I => \N__43954\
        );

    \I__9829\ : Span4Mux_v
    port map (
            O => \N__43957\,
            I => \N__43951\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43948\
        );

    \I__9827\ : Sp12to4
    port map (
            O => \N__43951\,
            I => \N__43942\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43942\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43939\
        );

    \I__9824\ : Span12Mux_h
    port map (
            O => \N__43942\,
            I => \N__43936\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43939\,
            I => buf_adcdata_vac_17
        );

    \I__9822\ : Odrv12
    port map (
            O => \N__43936\,
            I => buf_adcdata_vac_17
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__43931\,
            I => \n19_adj_1597_cascade_\
        );

    \I__9820\ : CascadeMux
    port map (
            O => \N__43928\,
            I => \n29_adj_1635_cascade_\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43925\,
            I => \N__43921\
        );

    \I__9818\ : CascadeMux
    port map (
            O => \N__43924\,
            I => \N__43917\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43921\,
            I => \N__43914\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43909\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43909\
        );

    \I__9814\ : Span4Mux_v
    port map (
            O => \N__43914\,
            I => \N__43904\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43909\,
            I => \N__43904\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__43904\,
            I => n16_adj_1623
        );

    \I__9811\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43896\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43891\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43891\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43896\,
            I => req_data_cnt_8
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43891\,
            I => req_data_cnt_8
        );

    \I__9806\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43883\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43883\,
            I => \N__43880\
        );

    \I__9804\ : Span4Mux_h
    port map (
            O => \N__43880\,
            I => \N__43875\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43872\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43869\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__43875\,
            I => n10534
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__43872\,
            I => n10534
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43869\,
            I => n10534
        );

    \I__9798\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43859\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43856\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43853\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__43853\,
            I => n20798
        );

    \I__9794\ : InMux
    port map (
            O => \N__43850\,
            I => \N__43847\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43847\,
            I => \N__43844\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__43844\,
            I => \N__43841\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__43841\,
            I => n22061
        );

    \I__9790\ : SRMux
    port map (
            O => \N__43838\,
            I => \N__43834\
        );

    \I__9789\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43831\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43828\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43825\
        );

    \I__9786\ : Odrv12
    port map (
            O => \N__43828\,
            I => n14730
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__43825\,
            I => n14730
        );

    \I__9784\ : ClkMux
    port map (
            O => \N__43820\,
            I => \N__43817\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43817\,
            I => \N__43810\
        );

    \I__9782\ : ClkMux
    port map (
            O => \N__43816\,
            I => \N__43807\
        );

    \I__9781\ : ClkMux
    port map (
            O => \N__43815\,
            I => \N__43801\
        );

    \I__9780\ : ClkMux
    port map (
            O => \N__43814\,
            I => \N__43798\
        );

    \I__9779\ : ClkMux
    port map (
            O => \N__43813\,
            I => \N__43795\
        );

    \I__9778\ : Span4Mux_v
    port map (
            O => \N__43810\,
            I => \N__43790\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43790\
        );

    \I__9776\ : ClkMux
    port map (
            O => \N__43806\,
            I => \N__43787\
        );

    \I__9775\ : ClkMux
    port map (
            O => \N__43805\,
            I => \N__43784\
        );

    \I__9774\ : ClkMux
    port map (
            O => \N__43804\,
            I => \N__43781\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43801\,
            I => \N__43776\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__43798\,
            I => \N__43773\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43795\,
            I => \N__43762\
        );

    \I__9770\ : Span4Mux_h
    port map (
            O => \N__43790\,
            I => \N__43762\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43787\,
            I => \N__43762\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__43784\,
            I => \N__43762\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43781\,
            I => \N__43762\
        );

    \I__9766\ : ClkMux
    port map (
            O => \N__43780\,
            I => \N__43755\
        );

    \I__9765\ : ClkMux
    port map (
            O => \N__43779\,
            I => \N__43752\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__43776\,
            I => \N__43749\
        );

    \I__9763\ : Span4Mux_v
    port map (
            O => \N__43773\,
            I => \N__43744\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__43762\,
            I => \N__43744\
        );

    \I__9761\ : ClkMux
    port map (
            O => \N__43761\,
            I => \N__43741\
        );

    \I__9760\ : ClkMux
    port map (
            O => \N__43760\,
            I => \N__43737\
        );

    \I__9759\ : ClkMux
    port map (
            O => \N__43759\,
            I => \N__43732\
        );

    \I__9758\ : ClkMux
    port map (
            O => \N__43758\,
            I => \N__43729\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43755\,
            I => \N__43726\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43752\,
            I => \N__43723\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__43749\,
            I => \N__43718\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__43744\,
            I => \N__43718\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43741\,
            I => \N__43715\
        );

    \I__9752\ : ClkMux
    port map (
            O => \N__43740\,
            I => \N__43712\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__43737\,
            I => \N__43709\
        );

    \I__9750\ : ClkMux
    port map (
            O => \N__43736\,
            I => \N__43706\
        );

    \I__9749\ : ClkMux
    port map (
            O => \N__43735\,
            I => \N__43703\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43732\,
            I => \N__43698\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43729\,
            I => \N__43698\
        );

    \I__9746\ : Span4Mux_h
    port map (
            O => \N__43726\,
            I => \N__43693\
        );

    \I__9745\ : Span4Mux_h
    port map (
            O => \N__43723\,
            I => \N__43693\
        );

    \I__9744\ : Span4Mux_h
    port map (
            O => \N__43718\,
            I => \N__43688\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__43715\,
            I => \N__43688\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43712\,
            I => \N__43685\
        );

    \I__9741\ : Span4Mux_h
    port map (
            O => \N__43709\,
            I => \N__43680\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__43706\,
            I => \N__43680\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__43703\,
            I => \N__43677\
        );

    \I__9738\ : Span4Mux_v
    port map (
            O => \N__43698\,
            I => \N__43674\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__43693\,
            I => \N__43671\
        );

    \I__9736\ : Sp12to4
    port map (
            O => \N__43688\,
            I => \N__43668\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__43685\,
            I => \N__43663\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__43680\,
            I => \N__43663\
        );

    \I__9733\ : Span4Mux_h
    port map (
            O => \N__43677\,
            I => \N__43660\
        );

    \I__9732\ : Span4Mux_h
    port map (
            O => \N__43674\,
            I => \N__43657\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__43671\,
            I => \N__43653\
        );

    \I__9730\ : Span12Mux_h
    port map (
            O => \N__43668\,
            I => \N__43650\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__43663\,
            I => \N__43647\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__43660\,
            I => \N__43644\
        );

    \I__9727\ : Span4Mux_h
    port map (
            O => \N__43657\,
            I => \N__43641\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43638\
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__43653\,
            I => \clk_RTD\
        );

    \I__9724\ : Odrv12
    port map (
            O => \N__43650\,
            I => \clk_RTD\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__43647\,
            I => \clk_RTD\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43644\,
            I => \clk_RTD\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__43641\,
            I => \clk_RTD\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43638\,
            I => \clk_RTD\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__43625\,
            I => \n22064_cascade_\
        );

    \I__9718\ : InMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__9716\ : Span4Mux_h
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9715\ : Span4Mux_h
    port map (
            O => \N__43613\,
            I => \N__43610\
        );

    \I__9714\ : Odrv4
    port map (
            O => \N__43610\,
            I => n16_adj_1519
        );

    \I__9713\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43604\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43604\,
            I => n22067
        );

    \I__9711\ : InMux
    port map (
            O => \N__43601\,
            I => \N__43597\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__43600\,
            I => \N__43594\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43591\
        );

    \I__9708\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43588\
        );

    \I__9707\ : Odrv12
    port map (
            O => \N__43591\,
            I => \buf_readRTD_5\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__43588\,
            I => \buf_readRTD_5\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43580\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__43580\,
            I => \N__43575\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43572\
        );

    \I__9702\ : CascadeMux
    port map (
            O => \N__43578\,
            I => \N__43569\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__43575\,
            I => \N__43566\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__43572\,
            I => \N__43563\
        );

    \I__9699\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43560\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__43566\,
            I => \N__43557\
        );

    \I__9697\ : Span12Mux_h
    port map (
            O => \N__43563\,
            I => \N__43554\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__43560\,
            I => buf_adcdata_iac_13
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__43557\,
            I => buf_adcdata_iac_13
        );

    \I__9694\ : Odrv12
    port map (
            O => \N__43554\,
            I => buf_adcdata_iac_13
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__43547\,
            I => \n22142_cascade_\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43541\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43541\,
            I => \N__43538\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__43538\,
            I => \N__43535\
        );

    \I__9689\ : Span4Mux_v
    port map (
            O => \N__43535\,
            I => \N__43532\
        );

    \I__9688\ : Odrv4
    port map (
            O => \N__43532\,
            I => n16_adj_1496
        );

    \I__9687\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43525\
        );

    \I__9686\ : CascadeMux
    port map (
            O => \N__43528\,
            I => \N__43521\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43525\,
            I => \N__43518\
        );

    \I__9684\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43515\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43521\,
            I => \N__43512\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__43518\,
            I => \N__43507\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43515\,
            I => \N__43507\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43512\,
            I => \acadc_skipCount_5\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__43507\,
            I => \acadc_skipCount_5\
        );

    \I__9678\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43499\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43499\,
            I => n22145
        );

    \I__9676\ : CascadeMux
    port map (
            O => \N__43496\,
            I => \n22133_cascade_\
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__43493\,
            I => \n30_adj_1499_cascade_\
        );

    \I__9674\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43486\
        );

    \I__9673\ : CascadeMux
    port map (
            O => \N__43489\,
            I => \N__43483\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__43486\,
            I => \N__43480\
        );

    \I__9671\ : InMux
    port map (
            O => \N__43483\,
            I => \N__43477\
        );

    \I__9670\ : Span4Mux_v
    port map (
            O => \N__43480\,
            I => \N__43474\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__43477\,
            I => data_idxvec_5
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__43474\,
            I => data_idxvec_5
        );

    \I__9667\ : CascadeMux
    port map (
            O => \N__43469\,
            I => \n26_adj_1498_cascade_\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43466\,
            I => \N__43463\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43463\,
            I => n22130
        );

    \I__9664\ : InMux
    port map (
            O => \N__43460\,
            I => \N__43455\
        );

    \I__9663\ : InMux
    port map (
            O => \N__43459\,
            I => \N__43452\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43458\,
            I => \N__43449\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__43455\,
            I => \N__43446\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__43452\,
            I => data_cntvec_8
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__43449\,
            I => data_cntvec_8
        );

    \I__9658\ : Odrv4
    port map (
            O => \N__43446\,
            I => data_cntvec_8
        );

    \I__9657\ : CascadeMux
    port map (
            O => \N__43439\,
            I => \N__43435\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43432\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43429\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__43432\,
            I => data_cntvec_13
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__43429\,
            I => data_cntvec_13
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__43424\,
            I => \n14545_cascade_\
        );

    \I__9651\ : CascadeMux
    port map (
            O => \N__43421\,
            I => \N__43417\
        );

    \I__9650\ : InMux
    port map (
            O => \N__43420\,
            I => \N__43414\
        );

    \I__9649\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43411\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43408\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43411\,
            I => data_idxvec_1
        );

    \I__9646\ : Odrv12
    port map (
            O => \N__43408\,
            I => data_idxvec_1
        );

    \I__9645\ : CascadeMux
    port map (
            O => \N__43403\,
            I => \n26_adj_1522_cascade_\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43400\,
            I => \N__43397\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43392\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43389\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43386\
        );

    \I__9640\ : Span4Mux_h
    port map (
            O => \N__43392\,
            I => \N__43381\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43381\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__43386\,
            I => \acadc_skipCount_1\
        );

    \I__9637\ : Odrv4
    port map (
            O => \N__43381\,
            I => \acadc_skipCount_1\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__43376\,
            I => \n22190_cascade_\
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__43373\,
            I => \n22193_cascade_\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__43370\,
            I => \n30_adj_1523_cascade_\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__43364\,
            I => \N__43361\
        );

    \I__9631\ : Span4Mux_v
    port map (
            O => \N__43361\,
            I => \N__43358\
        );

    \I__9630\ : Span4Mux_h
    port map (
            O => \N__43358\,
            I => \N__43355\
        );

    \I__9629\ : Odrv4
    port map (
            O => \N__43355\,
            I => n19_adj_1520
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__43352\,
            I => \N__43349\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43349\,
            I => \N__43346\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43346\,
            I => \N__43343\
        );

    \I__9625\ : Span4Mux_h
    port map (
            O => \N__43343\,
            I => \N__43340\
        );

    \I__9624\ : Sp12to4
    port map (
            O => \N__43340\,
            I => \N__43336\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43333\
        );

    \I__9622\ : Odrv12
    port map (
            O => \N__43336\,
            I => \buf_readRTD_1\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__43333\,
            I => \buf_readRTD_1\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43328\,
            I => \N__43325\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__43325\,
            I => \N__43322\
        );

    \I__9618\ : Span4Mux_h
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__43319\,
            I => comm_buf_5_2
        );

    \I__9616\ : InMux
    port map (
            O => \N__43316\,
            I => \N__43313\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43313\,
            I => \N__43310\
        );

    \I__9614\ : Odrv4
    port map (
            O => \N__43310\,
            I => comm_buf_4_2
        );

    \I__9613\ : InMux
    port map (
            O => \N__43307\,
            I => \N__43304\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__43304\,
            I => \N__43300\
        );

    \I__9611\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43297\
        );

    \I__9610\ : Span4Mux_v
    port map (
            O => \N__43300\,
            I => \N__43294\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43291\
        );

    \I__9608\ : Span4Mux_h
    port map (
            O => \N__43294\,
            I => \N__43288\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__43291\,
            I => comm_buf_6_2
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__43288\,
            I => comm_buf_6_2
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__43283\,
            I => \n4_adj_1593_cascade_\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43280\,
            I => \N__43277\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__43277\,
            I => n22049
        );

    \I__9602\ : CascadeMux
    port map (
            O => \N__43274\,
            I => \n20801_cascade_\
        );

    \I__9601\ : CascadeMux
    port map (
            O => \N__43271\,
            I => \N__43268\
        );

    \I__9600\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43265\,
            I => \N__43261\
        );

    \I__9598\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43258\
        );

    \I__9597\ : Odrv4
    port map (
            O => \N__43261\,
            I => n20596
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__43258\,
            I => n20596
        );

    \I__9595\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43250\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__43250\,
            I => \N__43247\
        );

    \I__9593\ : Span4Mux_v
    port map (
            O => \N__43247\,
            I => \N__43244\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__43244\,
            I => n21094
        );

    \I__9591\ : CascadeMux
    port map (
            O => \N__43241\,
            I => \n21092_cascade_\
        );

    \I__9590\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43235\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__43235\,
            I => n20_adj_1610
        );

    \I__9588\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__43229\,
            I => \N__43226\
        );

    \I__9586\ : Span4Mux_v
    port map (
            O => \N__43226\,
            I => \N__43223\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__43223\,
            I => n20883
        );

    \I__9584\ : CascadeMux
    port map (
            O => \N__43220\,
            I => \n20695_cascade_\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43214\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43214\,
            I => \N__43211\
        );

    \I__9581\ : Span4Mux_v
    port map (
            O => \N__43211\,
            I => \N__43208\
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__43208\,
            I => n20881
        );

    \I__9579\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__43202\,
            I => \N__43198\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43201\,
            I => \N__43195\
        );

    \I__9576\ : Span12Mux_v
    port map (
            O => \N__43198\,
            I => \N__43192\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__43195\,
            I => comm_buf_6_6
        );

    \I__9574\ : Odrv12
    port map (
            O => \N__43192\,
            I => comm_buf_6_6
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__43187\,
            I => \n21329_cascade_\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__43184\,
            I => \n21986_cascade_\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43178\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__43178\,
            I => n2_adj_1584
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__43175\,
            I => \N__43172\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43172\,
            I => \N__43169\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__43169\,
            I => \N__43165\
        );

    \I__9566\ : InMux
    port map (
            O => \N__43168\,
            I => \N__43162\
        );

    \I__9565\ : Span4Mux_v
    port map (
            O => \N__43165\,
            I => \N__43156\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43162\,
            I => \N__43156\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43161\,
            I => \N__43150\
        );

    \I__9562\ : Span4Mux_v
    port map (
            O => \N__43156\,
            I => \N__43146\
        );

    \I__9561\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43143\
        );

    \I__9560\ : InMux
    port map (
            O => \N__43154\,
            I => \N__43140\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43137\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__43150\,
            I => \N__43133\
        );

    \I__9557\ : InMux
    port map (
            O => \N__43149\,
            I => \N__43130\
        );

    \I__9556\ : Sp12to4
    port map (
            O => \N__43146\,
            I => \N__43125\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43125\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__43140\,
            I => \N__43122\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__43137\,
            I => \N__43119\
        );

    \I__9552\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43116\
        );

    \I__9551\ : Span4Mux_v
    port map (
            O => \N__43133\,
            I => \N__43111\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43130\,
            I => \N__43111\
        );

    \I__9549\ : Span12Mux_h
    port map (
            O => \N__43125\,
            I => \N__43108\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__43122\,
            I => \N__43103\
        );

    \I__9547\ : Span4Mux_h
    port map (
            O => \N__43119\,
            I => \N__43103\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__43116\,
            I => \N__43100\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__43111\,
            I => \N__43097\
        );

    \I__9544\ : Span12Mux_v
    port map (
            O => \N__43108\,
            I => \N__43094\
        );

    \I__9543\ : Span4Mux_v
    port map (
            O => \N__43103\,
            I => \N__43089\
        );

    \I__9542\ : Span4Mux_h
    port map (
            O => \N__43100\,
            I => \N__43089\
        );

    \I__9541\ : Span4Mux_h
    port map (
            O => \N__43097\,
            I => \N__43086\
        );

    \I__9540\ : Odrv12
    port map (
            O => \N__43094\,
            I => comm_buf_0_6
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__43089\,
            I => comm_buf_0_6
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__43086\,
            I => comm_buf_0_6
        );

    \I__9537\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__43076\,
            I => \N__43073\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__43073\,
            I => n1_adj_1583
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__43070\,
            I => \N__43067\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43064\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__43064\,
            I => \N__43060\
        );

    \I__9531\ : InMux
    port map (
            O => \N__43063\,
            I => \N__43056\
        );

    \I__9530\ : Span4Mux_v
    port map (
            O => \N__43060\,
            I => \N__43053\
        );

    \I__9529\ : InMux
    port map (
            O => \N__43059\,
            I => \N__43050\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__43056\,
            I => n20621
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__43053\,
            I => n20621
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__43050\,
            I => n20621
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__43043\,
            I => \n7_cascade_\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__43034\,
            I => \N__43031\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__43031\,
            I => \N__43028\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__43028\,
            I => comm_buf_2_2
        );

    \I__9519\ : CascadeMux
    port map (
            O => \N__43025\,
            I => \N__43022\
        );

    \I__9518\ : InMux
    port map (
            O => \N__43022\,
            I => \N__43019\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__43019\,
            I => \N__43016\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__43016\,
            I => \N__43013\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__43013\,
            I => comm_buf_3_2
        );

    \I__9514\ : CascadeMux
    port map (
            O => \N__43010\,
            I => \N__43006\
        );

    \I__9513\ : InMux
    port map (
            O => \N__43009\,
            I => \N__43000\
        );

    \I__9512\ : InMux
    port map (
            O => \N__43006\,
            I => \N__42997\
        );

    \I__9511\ : CascadeMux
    port map (
            O => \N__43005\,
            I => \N__42994\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__43004\,
            I => \N__42991\
        );

    \I__9509\ : CascadeMux
    port map (
            O => \N__43003\,
            I => \N__42988\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__43000\,
            I => \N__42982\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__42997\,
            I => \N__42982\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42979\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42976\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42988\,
            I => \N__42973\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42967\
        );

    \I__9502\ : Span4Mux_v
    port map (
            O => \N__42982\,
            I => \N__42962\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42979\,
            I => \N__42962\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42976\,
            I => \N__42959\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__42973\,
            I => \N__42956\
        );

    \I__9498\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42953\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42950\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42947\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42967\,
            I => \N__42944\
        );

    \I__9494\ : Span4Mux_v
    port map (
            O => \N__42962\,
            I => \N__42941\
        );

    \I__9493\ : Span4Mux_h
    port map (
            O => \N__42959\,
            I => \N__42936\
        );

    \I__9492\ : Span4Mux_v
    port map (
            O => \N__42956\,
            I => \N__42936\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__42953\,
            I => \N__42933\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__42950\,
            I => \N__42930\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42947\,
            I => \N__42923\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__42944\,
            I => \N__42923\
        );

    \I__9487\ : Span4Mux_h
    port map (
            O => \N__42941\,
            I => \N__42923\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__42936\,
            I => \N__42920\
        );

    \I__9485\ : Span4Mux_h
    port map (
            O => \N__42933\,
            I => \N__42917\
        );

    \I__9484\ : Span4Mux_h
    port map (
            O => \N__42930\,
            I => \N__42914\
        );

    \I__9483\ : Sp12to4
    port map (
            O => \N__42923\,
            I => \N__42911\
        );

    \I__9482\ : Span4Mux_h
    port map (
            O => \N__42920\,
            I => \N__42906\
        );

    \I__9481\ : Span4Mux_h
    port map (
            O => \N__42917\,
            I => \N__42906\
        );

    \I__9480\ : Span4Mux_h
    port map (
            O => \N__42914\,
            I => \N__42903\
        );

    \I__9479\ : Odrv12
    port map (
            O => \N__42911\,
            I => comm_buf_0_2
        );

    \I__9478\ : Odrv4
    port map (
            O => \N__42906\,
            I => comm_buf_0_2
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__42903\,
            I => comm_buf_0_2
        );

    \I__9476\ : CascadeMux
    port map (
            O => \N__42896\,
            I => \n22046_cascade_\
        );

    \I__9475\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42890\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42890\,
            I => \N__42887\
        );

    \I__9473\ : Span4Mux_h
    port map (
            O => \N__42887\,
            I => \N__42884\
        );

    \I__9472\ : Span4Mux_v
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__9471\ : Odrv4
    port map (
            O => \N__42881\,
            I => n30_adj_1529
        );

    \I__9470\ : InMux
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42872\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9467\ : Span4Mux_v
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__42866\,
            I => \N__42863\
        );

    \I__9465\ : Span4Mux_h
    port map (
            O => \N__42863\,
            I => \N__42860\
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__42860\,
            I => n22109
        );

    \I__9463\ : SRMux
    port map (
            O => \N__42857\,
            I => \N__42853\
        );

    \I__9462\ : SRMux
    port map (
            O => \N__42856\,
            I => \N__42848\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42853\,
            I => \N__42844\
        );

    \I__9460\ : SRMux
    port map (
            O => \N__42852\,
            I => \N__42841\
        );

    \I__9459\ : SRMux
    port map (
            O => \N__42851\,
            I => \N__42838\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__42848\,
            I => \N__42835\
        );

    \I__9457\ : SRMux
    port map (
            O => \N__42847\,
            I => \N__42832\
        );

    \I__9456\ : Span4Mux_v
    port map (
            O => \N__42844\,
            I => \N__42826\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42841\,
            I => \N__42826\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__42838\,
            I => \N__42823\
        );

    \I__9453\ : Span4Mux_h
    port map (
            O => \N__42835\,
            I => \N__42820\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42832\,
            I => \N__42817\
        );

    \I__9451\ : SRMux
    port map (
            O => \N__42831\,
            I => \N__42814\
        );

    \I__9450\ : Span4Mux_h
    port map (
            O => \N__42826\,
            I => \N__42811\
        );

    \I__9449\ : Span4Mux_h
    port map (
            O => \N__42823\,
            I => \N__42808\
        );

    \I__9448\ : Span4Mux_v
    port map (
            O => \N__42820\,
            I => \N__42803\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__42817\,
            I => \N__42803\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__42814\,
            I => \N__42800\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__42811\,
            I => n14766
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__42808\,
            I => n14766
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__42803\,
            I => n14766
        );

    \I__9442\ : Odrv12
    port map (
            O => \N__42800\,
            I => n14766
        );

    \I__9441\ : CascadeMux
    port map (
            O => \N__42791\,
            I => \n21199_cascade_\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__42788\,
            I => \n20681_cascade_\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42779\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42784\,
            I => \N__42773\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42773\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42770\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42779\,
            I => \N__42767\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42764\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42773\,
            I => \N__42761\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__42770\,
            I => \N__42758\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__42767\,
            I => \N__42755\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42764\,
            I => \N__42752\
        );

    \I__9429\ : Span4Mux_h
    port map (
            O => \N__42761\,
            I => \N__42749\
        );

    \I__9428\ : Span4Mux_h
    port map (
            O => \N__42758\,
            I => \N__42746\
        );

    \I__9427\ : Span4Mux_h
    port map (
            O => \N__42755\,
            I => \N__42741\
        );

    \I__9426\ : Span4Mux_h
    port map (
            O => \N__42752\,
            I => \N__42741\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__42749\,
            I => n20599
        );

    \I__9424\ : Odrv4
    port map (
            O => \N__42746\,
            I => n20599
        );

    \I__9423\ : Odrv4
    port map (
            O => \N__42741\,
            I => n20599
        );

    \I__9422\ : CascadeMux
    port map (
            O => \N__42734\,
            I => \n12108_cascade_\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42731\,
            I => \N__42728\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42728\,
            I => n4_adj_1616
        );

    \I__9419\ : CEMux
    port map (
            O => \N__42725\,
            I => \N__42718\
        );

    \I__9418\ : CEMux
    port map (
            O => \N__42724\,
            I => \N__42714\
        );

    \I__9417\ : CEMux
    port map (
            O => \N__42723\,
            I => \N__42711\
        );

    \I__9416\ : CEMux
    port map (
            O => \N__42722\,
            I => \N__42708\
        );

    \I__9415\ : CEMux
    port map (
            O => \N__42721\,
            I => \N__42705\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42718\,
            I => \N__42702\
        );

    \I__9413\ : CEMux
    port map (
            O => \N__42717\,
            I => \N__42699\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__42714\,
            I => \N__42696\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42711\,
            I => \N__42693\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__42708\,
            I => \N__42690\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__42705\,
            I => \N__42686\
        );

    \I__9408\ : Span12Mux_v
    port map (
            O => \N__42702\,
            I => \N__42683\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42699\,
            I => \N__42676\
        );

    \I__9406\ : Span4Mux_v
    port map (
            O => \N__42696\,
            I => \N__42676\
        );

    \I__9405\ : Span4Mux_v
    port map (
            O => \N__42693\,
            I => \N__42676\
        );

    \I__9404\ : Sp12to4
    port map (
            O => \N__42690\,
            I => \N__42673\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42689\,
            I => \N__42670\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__42686\,
            I => n11977
        );

    \I__9401\ : Odrv12
    port map (
            O => \N__42683\,
            I => n11977
        );

    \I__9400\ : Odrv4
    port map (
            O => \N__42676\,
            I => n11977
        );

    \I__9399\ : Odrv12
    port map (
            O => \N__42673\,
            I => n11977
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__42670\,
            I => n11977
        );

    \I__9397\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42656\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__9395\ : Span4Mux_h
    port map (
            O => \N__42653\,
            I => \N__42650\
        );

    \I__9394\ : Odrv4
    port map (
            O => \N__42650\,
            I => comm_buf_3_6
        );

    \I__9393\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42644\,
            I => \N__42641\
        );

    \I__9391\ : Odrv12
    port map (
            O => \N__42641\,
            I => comm_buf_2_6
        );

    \I__9390\ : InMux
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__42635\,
            I => \N__42632\
        );

    \I__9388\ : Odrv12
    port map (
            O => \N__42632\,
            I => buf_data_iac_22
        );

    \I__9387\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42626\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__42626\,
            I => \N__42623\
        );

    \I__9385\ : Span4Mux_v
    port map (
            O => \N__42623\,
            I => \N__42620\
        );

    \I__9384\ : Odrv4
    port map (
            O => \N__42620\,
            I => n21038
        );

    \I__9383\ : InMux
    port map (
            O => \N__42617\,
            I => \N__42614\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__42614\,
            I => \N__42611\
        );

    \I__9381\ : Span4Mux_v
    port map (
            O => \N__42611\,
            I => \N__42600\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42597\
        );

    \I__9379\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42582\
        );

    \I__9378\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42582\
        );

    \I__9377\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42582\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42582\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42582\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42582\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42582\
        );

    \I__9372\ : Odrv4
    port map (
            O => \N__42600\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42597\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__42582\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42568\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42574\,
            I => \N__42568\
        );

    \I__9367\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42565\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42568\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42565\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__9364\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42550\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42550\
        );

    \I__9362\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42550\
        );

    \I__9361\ : InMux
    port map (
            O => \N__42557\,
            I => \N__42547\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__42550\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__42547\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__9358\ : CascadeMux
    port map (
            O => \N__42542\,
            I => \N__42539\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42526\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42538\,
            I => \N__42526\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42537\,
            I => \N__42526\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42526\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42523\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42526\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__42523\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__9350\ : InMux
    port map (
            O => \N__42518\,
            I => n19507
        );

    \I__9349\ : InMux
    port map (
            O => \N__42515\,
            I => n19508
        );

    \I__9348\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42508\
        );

    \I__9347\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42505\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__42508\,
            I => clk_cnt_0
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__42505\,
            I => clk_cnt_0
        );

    \I__9344\ : InMux
    port map (
            O => \N__42500\,
            I => \N__42496\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42493\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__42496\,
            I => clk_cnt_4
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__42493\,
            I => clk_cnt_4
        );

    \I__9340\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42484\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42481\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42478\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__42481\,
            I => clk_cnt_1
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__42478\,
            I => clk_cnt_1
        );

    \I__9335\ : InMux
    port map (
            O => \N__42473\,
            I => \N__42469\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42466\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__42469\,
            I => clk_cnt_3
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__42466\,
            I => clk_cnt_3
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__42461\,
            I => \n6_cascade_\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42454\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42451\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42448\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__42451\,
            I => clk_cnt_2
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__42448\,
            I => clk_cnt_2
        );

    \I__9325\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42440\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42440\,
            I => \N__42435\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__42439\,
            I => \N__42432\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__42438\,
            I => \N__42429\
        );

    \I__9321\ : Span4Mux_h
    port map (
            O => \N__42435\,
            I => \N__42426\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42421\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42421\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__42426\,
            I => \acadc_skipCount_11\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__42421\,
            I => \acadc_skipCount_11\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42412\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42415\,
            I => \N__42409\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__42412\,
            I => dds0_mclkcnt_3
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42409\,
            I => dds0_mclkcnt_3
        );

    \I__9312\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42400\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42397\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__42400\,
            I => dds0_mclkcnt_5
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__42397\,
            I => dds0_mclkcnt_5
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__42392\,
            I => \N__42388\
        );

    \I__9307\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42385\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42388\,
            I => \N__42382\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42385\,
            I => dds0_mclkcnt_1
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42382\,
            I => dds0_mclkcnt_1
        );

    \I__9303\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42373\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42370\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__42373\,
            I => dds0_mclkcnt_4
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42370\,
            I => dds0_mclkcnt_4
        );

    \I__9299\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42361\
        );

    \I__9298\ : InMux
    port map (
            O => \N__42364\,
            I => \N__42358\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__42361\,
            I => dds0_mclkcnt_2
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42358\,
            I => dds0_mclkcnt_2
        );

    \I__9295\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42349\
        );

    \I__9294\ : InMux
    port map (
            O => \N__42352\,
            I => \N__42346\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__42349\,
            I => dds0_mclkcnt_0
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__42346\,
            I => dds0_mclkcnt_0
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__42341\,
            I => \n12_cascade_\
        );

    \I__9290\ : InMux
    port map (
            O => \N__42338\,
            I => \N__42334\
        );

    \I__9289\ : InMux
    port map (
            O => \N__42337\,
            I => \N__42331\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__42334\,
            I => dds0_mclkcnt_7
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42331\,
            I => dds0_mclkcnt_7
        );

    \I__9286\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42323\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__42323\,
            I => n20543
        );

    \I__9284\ : CascadeMux
    port map (
            O => \N__42320\,
            I => \n20543_cascade_\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42313\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42310\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42313\,
            I => dds0_mclkcnt_6
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42310\,
            I => dds0_mclkcnt_6
        );

    \I__9279\ : CascadeMux
    port map (
            O => \N__42305\,
            I => \n8_adj_1559_cascade_\
        );

    \I__9278\ : CascadeMux
    port map (
            O => \N__42302\,
            I => \N__42299\
        );

    \I__9277\ : CascadeBuf
    port map (
            O => \N__42299\,
            I => \N__42296\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \N__42293\
        );

    \I__9275\ : CascadeBuf
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__42290\,
            I => \N__42287\
        );

    \I__9273\ : CascadeBuf
    port map (
            O => \N__42287\,
            I => \N__42284\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__9271\ : CascadeBuf
    port map (
            O => \N__42281\,
            I => \N__42278\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__42278\,
            I => \N__42275\
        );

    \I__9269\ : CascadeBuf
    port map (
            O => \N__42275\,
            I => \N__42272\
        );

    \I__9268\ : CascadeMux
    port map (
            O => \N__42272\,
            I => \N__42269\
        );

    \I__9267\ : CascadeBuf
    port map (
            O => \N__42269\,
            I => \N__42266\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__42266\,
            I => \N__42263\
        );

    \I__9265\ : CascadeBuf
    port map (
            O => \N__42263\,
            I => \N__42260\
        );

    \I__9264\ : CascadeMux
    port map (
            O => \N__42260\,
            I => \N__42256\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__42259\,
            I => \N__42253\
        );

    \I__9262\ : CascadeBuf
    port map (
            O => \N__42256\,
            I => \N__42250\
        );

    \I__9261\ : CascadeBuf
    port map (
            O => \N__42253\,
            I => \N__42247\
        );

    \I__9260\ : CascadeMux
    port map (
            O => \N__42250\,
            I => \N__42244\
        );

    \I__9259\ : CascadeMux
    port map (
            O => \N__42247\,
            I => \N__42241\
        );

    \I__9258\ : CascadeBuf
    port map (
            O => \N__42244\,
            I => \N__42238\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42235\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__42238\,
            I => \N__42232\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__42235\,
            I => \N__42229\
        );

    \I__9254\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42226\
        );

    \I__9253\ : Span12Mux_h
    port map (
            O => \N__42229\,
            I => \N__42223\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__42226\,
            I => \N__42220\
        );

    \I__9251\ : Span12Mux_v
    port map (
            O => \N__42223\,
            I => \N__42215\
        );

    \I__9250\ : Span12Mux_s11_v
    port map (
            O => \N__42220\,
            I => \N__42215\
        );

    \I__9249\ : Odrv12
    port map (
            O => \N__42215\,
            I => \data_index_9_N_216_6\
        );

    \I__9248\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42209\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42206\
        );

    \I__9246\ : Span4Mux_v
    port map (
            O => \N__42206\,
            I => \N__42203\
        );

    \I__9245\ : Odrv4
    port map (
            O => \N__42203\,
            I => n8_adj_1567
        );

    \I__9244\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42196\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42193\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42196\,
            I => \N__42190\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42193\,
            I => \N__42187\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__42190\,
            I => \N__42182\
        );

    \I__9239\ : Span4Mux_h
    port map (
            O => \N__42187\,
            I => \N__42182\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__42182\,
            I => \N__42179\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__42179\,
            I => n7_adj_1566
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__42176\,
            I => \N__42173\
        );

    \I__9235\ : CascadeBuf
    port map (
            O => \N__42173\,
            I => \N__42170\
        );

    \I__9234\ : CascadeMux
    port map (
            O => \N__42170\,
            I => \N__42167\
        );

    \I__9233\ : CascadeBuf
    port map (
            O => \N__42167\,
            I => \N__42164\
        );

    \I__9232\ : CascadeMux
    port map (
            O => \N__42164\,
            I => \N__42161\
        );

    \I__9231\ : CascadeBuf
    port map (
            O => \N__42161\,
            I => \N__42158\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__42158\,
            I => \N__42155\
        );

    \I__9229\ : CascadeBuf
    port map (
            O => \N__42155\,
            I => \N__42152\
        );

    \I__9228\ : CascadeMux
    port map (
            O => \N__42152\,
            I => \N__42149\
        );

    \I__9227\ : CascadeBuf
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__9226\ : CascadeMux
    port map (
            O => \N__42146\,
            I => \N__42143\
        );

    \I__9225\ : CascadeBuf
    port map (
            O => \N__42143\,
            I => \N__42140\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__42140\,
            I => \N__42137\
        );

    \I__9223\ : CascadeBuf
    port map (
            O => \N__42137\,
            I => \N__42134\
        );

    \I__9222\ : CascadeMux
    port map (
            O => \N__42134\,
            I => \N__42131\
        );

    \I__9221\ : CascadeBuf
    port map (
            O => \N__42131\,
            I => \N__42127\
        );

    \I__9220\ : CascadeMux
    port map (
            O => \N__42130\,
            I => \N__42124\
        );

    \I__9219\ : CascadeMux
    port map (
            O => \N__42127\,
            I => \N__42121\
        );

    \I__9218\ : CascadeBuf
    port map (
            O => \N__42124\,
            I => \N__42118\
        );

    \I__9217\ : CascadeBuf
    port map (
            O => \N__42121\,
            I => \N__42115\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__42118\,
            I => \N__42112\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__42115\,
            I => \N__42109\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42112\,
            I => \N__42106\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42103\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42100\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__42103\,
            I => \N__42097\
        );

    \I__9210\ : Span12Mux_s11_h
    port map (
            O => \N__42100\,
            I => \N__42094\
        );

    \I__9209\ : Span4Mux_h
    port map (
            O => \N__42097\,
            I => \N__42091\
        );

    \I__9208\ : Span12Mux_v
    port map (
            O => \N__42094\,
            I => \N__42088\
        );

    \I__9207\ : Span4Mux_v
    port map (
            O => \N__42091\,
            I => \N__42085\
        );

    \I__9206\ : Odrv12
    port map (
            O => \N__42088\,
            I => \data_index_9_N_216_1\
        );

    \I__9205\ : Odrv4
    port map (
            O => \N__42085\,
            I => \data_index_9_N_216_1\
        );

    \I__9204\ : InMux
    port map (
            O => \N__42080\,
            I => \N__42076\
        );

    \I__9203\ : InMux
    port map (
            O => \N__42079\,
            I => \N__42073\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__42076\,
            I => data_cntvec_12
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__42073\,
            I => data_cntvec_12
        );

    \I__9200\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42065\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__42065\,
            I => \N__42062\
        );

    \I__9198\ : Span4Mux_h
    port map (
            O => \N__42062\,
            I => \N__42057\
        );

    \I__9197\ : InMux
    port map (
            O => \N__42061\,
            I => \N__42054\
        );

    \I__9196\ : InMux
    port map (
            O => \N__42060\,
            I => \N__42051\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__42057\,
            I => \N__42048\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__42054\,
            I => data_cntvec_10
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__42051\,
            I => data_cntvec_10
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__42048\,
            I => data_cntvec_10
        );

    \I__9191\ : InMux
    port map (
            O => \N__42041\,
            I => \N__42036\
        );

    \I__9190\ : CascadeMux
    port map (
            O => \N__42040\,
            I => \N__42033\
        );

    \I__9189\ : InMux
    port map (
            O => \N__42039\,
            I => \N__42030\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__42036\,
            I => \N__42027\
        );

    \I__9187\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42024\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__42030\,
            I => req_data_cnt_12
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__42027\,
            I => req_data_cnt_12
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__42024\,
            I => req_data_cnt_12
        );

    \I__9183\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42014\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__42014\,
            I => \N__42010\
        );

    \I__9181\ : InMux
    port map (
            O => \N__42013\,
            I => \N__42006\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__42010\,
            I => \N__42003\
        );

    \I__9179\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42000\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__42006\,
            I => req_data_cnt_10
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__42003\,
            I => req_data_cnt_10
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__42000\,
            I => req_data_cnt_10
        );

    \I__9175\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41990\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41990\,
            I => n8_adj_1559
        );

    \I__9173\ : CascadeMux
    port map (
            O => \N__41987\,
            I => \N__41984\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41978\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41978\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41978\,
            I => \N__41975\
        );

    \I__9169\ : Span4Mux_v
    port map (
            O => \N__41975\,
            I => \N__41972\
        );

    \I__9168\ : Span4Mux_v
    port map (
            O => \N__41972\,
            I => \N__41969\
        );

    \I__9167\ : Span4Mux_h
    port map (
            O => \N__41969\,
            I => \N__41966\
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__41966\,
            I => n7_adj_1558
        );

    \I__9165\ : InMux
    port map (
            O => \N__41963\,
            I => \N__41959\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41962\,
            I => \N__41956\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41959\,
            I => \N__41953\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41956\,
            I => \N__41950\
        );

    \I__9161\ : Span4Mux_h
    port map (
            O => \N__41953\,
            I => \N__41946\
        );

    \I__9160\ : Span4Mux_h
    port map (
            O => \N__41950\,
            I => \N__41943\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41940\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__41946\,
            I => \N__41935\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__41943\,
            I => \N__41935\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__41940\,
            I => data_index_6
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__41935\,
            I => data_index_6
        );

    \I__9154\ : SRMux
    port map (
            O => \N__41930\,
            I => \N__41927\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__41927\,
            I => \N__41924\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__41924\,
            I => \N__41921\
        );

    \I__9151\ : Span4Mux_v
    port map (
            O => \N__41921\,
            I => \N__41918\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__41918\,
            I => \comm_spi.data_tx_7__N_771\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41915\,
            I => \bfn_15_16_0_\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41912\,
            I => n19505
        );

    \I__9147\ : InMux
    port map (
            O => \N__41909\,
            I => n19506
        );

    \I__9146\ : InMux
    port map (
            O => \N__41906\,
            I => n19363
        );

    \I__9145\ : InMux
    port map (
            O => \N__41903\,
            I => n19364
        );

    \I__9144\ : InMux
    port map (
            O => \N__41900\,
            I => n19365
        );

    \I__9143\ : InMux
    port map (
            O => \N__41897\,
            I => n19366
        );

    \I__9142\ : InMux
    port map (
            O => \N__41894\,
            I => n19367
        );

    \I__9141\ : InMux
    port map (
            O => \N__41891\,
            I => n19368
        );

    \I__9140\ : CEMux
    port map (
            O => \N__41888\,
            I => \N__41882\
        );

    \I__9139\ : CEMux
    port map (
            O => \N__41887\,
            I => \N__41879\
        );

    \I__9138\ : CEMux
    port map (
            O => \N__41886\,
            I => \N__41876\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41872\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41882\,
            I => \N__41869\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41879\,
            I => \N__41866\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41876\,
            I => \N__41863\
        );

    \I__9133\ : CEMux
    port map (
            O => \N__41875\,
            I => \N__41860\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__41872\,
            I => \N__41857\
        );

    \I__9131\ : Span4Mux_v
    port map (
            O => \N__41869\,
            I => \N__41848\
        );

    \I__9130\ : Span4Mux_v
    port map (
            O => \N__41866\,
            I => \N__41848\
        );

    \I__9129\ : Span4Mux_v
    port map (
            O => \N__41863\,
            I => \N__41848\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41848\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__41857\,
            I => \N__41845\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__41848\,
            I => n13473
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__41845\,
            I => n13473
        );

    \I__9124\ : SRMux
    port map (
            O => \N__41840\,
            I => \N__41836\
        );

    \I__9123\ : SRMux
    port map (
            O => \N__41839\,
            I => \N__41833\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41836\,
            I => \N__41829\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41833\,
            I => \N__41825\
        );

    \I__9120\ : SRMux
    port map (
            O => \N__41832\,
            I => \N__41822\
        );

    \I__9119\ : Span4Mux_h
    port map (
            O => \N__41829\,
            I => \N__41819\
        );

    \I__9118\ : SRMux
    port map (
            O => \N__41828\,
            I => \N__41816\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__41825\,
            I => \N__41811\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41822\,
            I => \N__41811\
        );

    \I__9115\ : Sp12to4
    port map (
            O => \N__41819\,
            I => \N__41806\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41816\,
            I => \N__41806\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__41811\,
            I => \N__41803\
        );

    \I__9112\ : Odrv12
    port map (
            O => \N__41806\,
            I => n14663
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__41803\,
            I => n14663
        );

    \I__9110\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41794\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41791\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__41794\,
            I => data_cntvec_14
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41791\,
            I => data_cntvec_14
        );

    \I__9106\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41781\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41778\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41775\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__41781\,
            I => \N__41772\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41778\,
            I => data_cntvec_11
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__41775\,
            I => data_cntvec_11
        );

    \I__9100\ : Odrv12
    port map (
            O => \N__41772\,
            I => data_cntvec_11
        );

    \I__9099\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41758\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41758\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41755\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__41758\,
            I => req_data_cnt_14
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41755\,
            I => req_data_cnt_14
        );

    \I__9094\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41743\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41740\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41748\,
            I => \N__41737\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41747\,
            I => \N__41734\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41731\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41743\,
            I => \N__41725\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41722\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41737\,
            I => \N__41715\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41734\,
            I => \N__41715\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__41731\,
            I => \N__41715\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41710\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41729\,
            I => \N__41710\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41728\,
            I => \N__41705\
        );

    \I__9081\ : Span4Mux_h
    port map (
            O => \N__41725\,
            I => \N__41696\
        );

    \I__9080\ : Span4Mux_h
    port map (
            O => \N__41722\,
            I => \N__41696\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__41715\,
            I => \N__41696\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41710\,
            I => \N__41696\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41709\,
            I => \N__41691\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41691\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41705\,
            I => n8828
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__41696\,
            I => n8828
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__41691\,
            I => n8828
        );

    \I__9072\ : InMux
    port map (
            O => \N__41684\,
            I => n19354
        );

    \I__9071\ : InMux
    port map (
            O => \N__41681\,
            I => n19355
        );

    \I__9070\ : InMux
    port map (
            O => \N__41678\,
            I => n19356
        );

    \I__9069\ : InMux
    port map (
            O => \N__41675\,
            I => n19357
        );

    \I__9068\ : InMux
    port map (
            O => \N__41672\,
            I => n19358
        );

    \I__9067\ : InMux
    port map (
            O => \N__41669\,
            I => n19359
        );

    \I__9066\ : InMux
    port map (
            O => \N__41666\,
            I => n19360
        );

    \I__9065\ : InMux
    port map (
            O => \N__41663\,
            I => \bfn_15_14_0_\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41660\,
            I => n19362
        );

    \I__9063\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41653\
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__41656\,
            I => \N__41650\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41653\,
            I => \N__41647\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41643\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__41647\,
            I => \N__41640\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41637\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__41643\,
            I => \acadc_skipCount_8\
        );

    \I__9056\ : Odrv4
    port map (
            O => \N__41640\,
            I => \acadc_skipCount_8\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41637\,
            I => \acadc_skipCount_8\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41627\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__41627\,
            I => \N__41620\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41615\
        );

    \I__9051\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41615\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41612\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41609\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__41620\,
            I => \N__41606\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__41615\,
            I => \N__41603\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41600\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__41609\,
            I => eis_start
        );

    \I__9044\ : Odrv4
    port map (
            O => \N__41606\,
            I => eis_start
        );

    \I__9043\ : Odrv4
    port map (
            O => \N__41603\,
            I => eis_start
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__41600\,
            I => eis_start
        );

    \I__9041\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41588\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__41588\,
            I => n21992
        );

    \I__9039\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41581\
        );

    \I__9038\ : CascadeMux
    port map (
            O => \N__41584\,
            I => \N__41578\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41575\
        );

    \I__9036\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41572\
        );

    \I__9035\ : Span4Mux_h
    port map (
            O => \N__41575\,
            I => \N__41569\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41572\,
            I => data_idxvec_8
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__41569\,
            I => data_idxvec_8
        );

    \I__9032\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41561\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41561\,
            I => \N__41558\
        );

    \I__9030\ : Odrv12
    port map (
            O => \N__41558\,
            I => buf_data_iac_16
        );

    \I__9029\ : CascadeMux
    port map (
            O => \N__41555\,
            I => \n20917_cascade_\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41552\,
            I => \N__41549\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41549\,
            I => n21995
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__41546\,
            I => \n20919_cascade_\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41540\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41537\
        );

    \I__9023\ : Span12Mux_h
    port map (
            O => \N__41537\,
            I => \N__41534\
        );

    \I__9022\ : Odrv12
    port map (
            O => \N__41534\,
            I => n22043
        );

    \I__9021\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41528\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41528\,
            I => \N__41525\
        );

    \I__9019\ : Span4Mux_v
    port map (
            O => \N__41525\,
            I => \N__41522\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__41522\,
            I => \N__41519\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__41519\,
            I => n22019
        );

    \I__9016\ : CascadeMux
    port map (
            O => \N__41516\,
            I => \n22220_cascade_\
        );

    \I__9015\ : CascadeMux
    port map (
            O => \N__41513\,
            I => \n22223_cascade_\
        );

    \I__9014\ : CascadeMux
    port map (
            O => \N__41510\,
            I => \N__41507\
        );

    \I__9013\ : InMux
    port map (
            O => \N__41507\,
            I => \N__41501\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41501\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41501\,
            I => \N__41495\
        );

    \I__9010\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41490\
        );

    \I__9009\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41487\
        );

    \I__9008\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41484\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__41495\,
            I => \N__41481\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41478\
        );

    \I__9005\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41475\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41472\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__41487\,
            I => \N__41469\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__41484\,
            I => \N__41466\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__41481\,
            I => \N__41461\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41478\,
            I => \N__41461\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41475\,
            I => \N__41456\
        );

    \I__8998\ : Span4Mux_v
    port map (
            O => \N__41472\,
            I => \N__41456\
        );

    \I__8997\ : Span4Mux_h
    port map (
            O => \N__41469\,
            I => \N__41451\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__41466\,
            I => \N__41451\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__41461\,
            I => \N__41444\
        );

    \I__8994\ : Span4Mux_v
    port map (
            O => \N__41456\,
            I => \N__41444\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__41451\,
            I => \N__41444\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__41444\,
            I => comm_buf_0_0
        );

    \I__8991\ : CascadeMux
    port map (
            O => \N__41441\,
            I => \N__41438\
        );

    \I__8990\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41434\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41429\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41434\,
            I => \N__41426\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41423\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41420\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41415\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__41426\,
            I => \N__41412\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__41423\,
            I => \N__41407\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41407\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41419\,
            I => \N__41402\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41418\,
            I => \N__41402\
        );

    \I__8979\ : Span4Mux_v
    port map (
            O => \N__41415\,
            I => \N__41395\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__41412\,
            I => \N__41395\
        );

    \I__8977\ : Span4Mux_v
    port map (
            O => \N__41407\,
            I => \N__41395\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__41402\,
            I => \iac_raw_buf_N_737\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__41395\,
            I => \iac_raw_buf_N_737\
        );

    \I__8974\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41383\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41389\,
            I => \N__41383\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41388\,
            I => \N__41379\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41376\
        );

    \I__8970\ : CascadeMux
    port map (
            O => \N__41382\,
            I => \N__41372\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41379\,
            I => \N__41367\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__41376\,
            I => \N__41364\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41361\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41358\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41353\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41353\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__41367\,
            I => \N__41348\
        );

    \I__8962\ : Span4Mux_h
    port map (
            O => \N__41364\,
            I => \N__41348\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41361\,
            I => n12397
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41358\,
            I => n12397
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__41353\,
            I => n12397
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__41348\,
            I => n12397
        );

    \I__8957\ : IoInMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__8955\ : Span4Mux_s2_h
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__8954\ : Span4Mux_h
    port map (
            O => \N__41330\,
            I => \N__41327\
        );

    \I__8953\ : Sp12to4
    port map (
            O => \N__41327\,
            I => \N__41324\
        );

    \I__8952\ : Span12Mux_s10_v
    port map (
            O => \N__41324\,
            I => \N__41319\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41316\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41313\
        );

    \I__8949\ : Span12Mux_h
    port map (
            O => \N__41319\,
            I => \N__41308\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__41316\,
            I => \N__41308\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__41313\,
            I => \VAC_OSR0\
        );

    \I__8946\ : Odrv12
    port map (
            O => \N__41308\,
            I => \VAC_OSR0\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41300\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__41300\,
            I => \N__41297\
        );

    \I__8943\ : Span4Mux_v
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__8942\ : Odrv4
    port map (
            O => \N__41294\,
            I => n21046
        );

    \I__8941\ : InMux
    port map (
            O => \N__41291\,
            I => \N__41288\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__8939\ : Span4Mux_h
    port map (
            O => \N__41285\,
            I => \N__41280\
        );

    \I__8938\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41275\
        );

    \I__8937\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41275\
        );

    \I__8936\ : Odrv4
    port map (
            O => \N__41280\,
            I => \acadc_skipCount_0\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__41275\,
            I => \acadc_skipCount_0\
        );

    \I__8934\ : InMux
    port map (
            O => \N__41270\,
            I => \N__41267\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41267\,
            I => \N__41264\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__41264\,
            I => \N__41261\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__41261\,
            I => n19_adj_1487
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__41258\,
            I => \N__41255\
        );

    \I__8929\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41252\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__41252\,
            I => \N__41248\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__41251\,
            I => \N__41245\
        );

    \I__8926\ : Span12Mux_h
    port map (
            O => \N__41248\,
            I => \N__41242\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41239\
        );

    \I__8924\ : Odrv12
    port map (
            O => \N__41242\,
            I => \buf_readRTD_0\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__41239\,
            I => \buf_readRTD_0\
        );

    \I__8922\ : CascadeMux
    port map (
            O => \N__41234\,
            I => \N__41230\
        );

    \I__8921\ : InMux
    port map (
            O => \N__41233\,
            I => \N__41227\
        );

    \I__8920\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41224\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41221\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41224\,
            I => data_idxvec_0
        );

    \I__8917\ : Odrv12
    port map (
            O => \N__41221\,
            I => data_idxvec_0
        );

    \I__8916\ : InMux
    port map (
            O => \N__41216\,
            I => \N__41213\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__41213\,
            I => \N__41210\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__41210\,
            I => n20973
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__41207\,
            I => \n26_cascade_\
        );

    \I__8912\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41201\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__41201\,
            I => n21998
        );

    \I__8910\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41195\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__41195\,
            I => \N__41192\
        );

    \I__8908\ : Span4Mux_h
    port map (
            O => \N__41192\,
            I => \N__41189\
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__41189\,
            I => n16_adj_1488
        );

    \I__8906\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__41183\,
            I => n22004
        );

    \I__8904\ : CascadeMux
    port map (
            O => \N__41180\,
            I => \n22007_cascade_\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__41174\,
            I => n22001
        );

    \I__8901\ : CascadeMux
    port map (
            O => \N__41171\,
            I => \n30_adj_1486_cascade_\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__41168\,
            I => \N__41164\
        );

    \I__8899\ : CascadeMux
    port map (
            O => \N__41167\,
            I => \N__41159\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41150\
        );

    \I__8897\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41150\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41150\
        );

    \I__8895\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41147\
        );

    \I__8894\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41144\
        );

    \I__8893\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41141\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41138\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41147\,
            I => \N__41133\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41144\,
            I => \N__41133\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41141\,
            I => \N__41130\
        );

    \I__8888\ : Span4Mux_h
    port map (
            O => \N__41138\,
            I => \N__41127\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__41133\,
            I => \N__41124\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__41130\,
            I => \N__41121\
        );

    \I__8885\ : Span4Mux_h
    port map (
            O => \N__41127\,
            I => \N__41118\
        );

    \I__8884\ : Span4Mux_v
    port map (
            O => \N__41124\,
            I => \N__41115\
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__41121\,
            I => comm_buf_1_0
        );

    \I__8882\ : Odrv4
    port map (
            O => \N__41118\,
            I => comm_buf_1_0
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__41115\,
            I => comm_buf_1_0
        );

    \I__8880\ : CascadeMux
    port map (
            O => \N__41108\,
            I => \n12242_cascade_\
        );

    \I__8879\ : CascadeMux
    port map (
            O => \N__41105\,
            I => \n20599_cascade_\
        );

    \I__8878\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41099\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__41099\,
            I => \N__41096\
        );

    \I__8876\ : Odrv12
    port map (
            O => \N__41096\,
            I => n5
        );

    \I__8875\ : IoInMux
    port map (
            O => \N__41093\,
            I => \N__41090\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__41090\,
            I => \N__41087\
        );

    \I__8873\ : IoSpan4Mux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__8872\ : Span4Mux_s3_v
    port map (
            O => \N__41084\,
            I => \N__41081\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__41081\,
            I => \N__41078\
        );

    \I__8870\ : Sp12to4
    port map (
            O => \N__41078\,
            I => \N__41074\
        );

    \I__8869\ : InMux
    port map (
            O => \N__41077\,
            I => \N__41070\
        );

    \I__8868\ : Span12Mux_h
    port map (
            O => \N__41074\,
            I => \N__41067\
        );

    \I__8867\ : InMux
    port map (
            O => \N__41073\,
            I => \N__41064\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__41070\,
            I => \N__41061\
        );

    \I__8865\ : Odrv12
    port map (
            O => \N__41067\,
            I => \IAC_FLT1\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__41064\,
            I => \IAC_FLT1\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__41061\,
            I => \IAC_FLT1\
        );

    \I__8862\ : CascadeMux
    port map (
            O => \N__41054\,
            I => \N__41046\
        );

    \I__8861\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41042\
        );

    \I__8860\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41037\
        );

    \I__8859\ : InMux
    port map (
            O => \N__41051\,
            I => \N__41037\
        );

    \I__8858\ : CascadeMux
    port map (
            O => \N__41050\,
            I => \N__41032\
        );

    \I__8857\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41027\
        );

    \I__8856\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41027\
        );

    \I__8855\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41024\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41017\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__41037\,
            I => \N__41014\
        );

    \I__8852\ : InMux
    port map (
            O => \N__41036\,
            I => \N__41011\
        );

    \I__8851\ : InMux
    port map (
            O => \N__41035\,
            I => \N__41006\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41006\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__41027\,
            I => \N__41003\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__41024\,
            I => \N__41000\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41023\,
            I => \N__40997\
        );

    \I__8846\ : InMux
    port map (
            O => \N__41022\,
            I => \N__40994\
        );

    \I__8845\ : InMux
    port map (
            O => \N__41021\,
            I => \N__40991\
        );

    \I__8844\ : InMux
    port map (
            O => \N__41020\,
            I => \N__40988\
        );

    \I__8843\ : Span4Mux_h
    port map (
            O => \N__41017\,
            I => \N__40985\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__41014\,
            I => \N__40982\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__41011\,
            I => \N__40973\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__41006\,
            I => \N__40973\
        );

    \I__8839\ : Span4Mux_h
    port map (
            O => \N__41003\,
            I => \N__40973\
        );

    \I__8838\ : Span4Mux_h
    port map (
            O => \N__41000\,
            I => \N__40973\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40997\,
            I => eis_state_1
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40994\,
            I => eis_state_1
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40991\,
            I => eis_state_1
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__40988\,
            I => eis_state_1
        );

    \I__8833\ : Odrv4
    port map (
            O => \N__40985\,
            I => eis_state_1
        );

    \I__8832\ : Odrv4
    port map (
            O => \N__40982\,
            I => eis_state_1
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__40973\,
            I => eis_state_1
        );

    \I__8830\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40955\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40952\
        );

    \I__8828\ : Span12Mux_h
    port map (
            O => \N__40952\,
            I => \N__40949\
        );

    \I__8827\ : Odrv12
    port map (
            O => \N__40949\,
            I => buf_data_iac_8
        );

    \I__8826\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40942\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__40945\,
            I => \N__40939\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40936\
        );

    \I__8823\ : InMux
    port map (
            O => \N__40939\,
            I => \N__40933\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__40936\,
            I => \N__40930\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40933\,
            I => data_idxvec_12
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__40930\,
            I => data_idxvec_12
        );

    \I__8819\ : CascadeMux
    port map (
            O => \N__40925\,
            I => \N__40922\
        );

    \I__8818\ : InMux
    port map (
            O => \N__40922\,
            I => \N__40919\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__40919\,
            I => \N__40916\
        );

    \I__8816\ : Odrv12
    port map (
            O => \N__40916\,
            I => n20983
        );

    \I__8815\ : InMux
    port map (
            O => \N__40913\,
            I => \N__40910\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40910\,
            I => \N__40906\
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__40909\,
            I => \N__40903\
        );

    \I__8812\ : Span4Mux_h
    port map (
            O => \N__40906\,
            I => \N__40900\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40897\
        );

    \I__8810\ : Span4Mux_v
    port map (
            O => \N__40900\,
            I => \N__40894\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__40897\,
            I => \N__40890\
        );

    \I__8808\ : Span4Mux_h
    port map (
            O => \N__40894\,
            I => \N__40887\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40884\
        );

    \I__8806\ : Span12Mux_v
    port map (
            O => \N__40890\,
            I => \N__40881\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__40887\,
            I => \N__40878\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40884\,
            I => buf_adcdata_iac_19
        );

    \I__8803\ : Odrv12
    port map (
            O => \N__40881\,
            I => buf_adcdata_iac_19
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__40878\,
            I => buf_adcdata_iac_19
        );

    \I__8801\ : InMux
    port map (
            O => \N__40871\,
            I => \N__40868\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__40868\,
            I => n22082
        );

    \I__8799\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40861\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__40864\,
            I => \N__40858\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40855\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40858\,
            I => \N__40852\
        );

    \I__8795\ : Span4Mux_h
    port map (
            O => \N__40855\,
            I => \N__40849\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40852\,
            I => data_idxvec_11
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__40849\,
            I => data_idxvec_11
        );

    \I__8792\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40841\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__40841\,
            I => \N__40838\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__40838\,
            I => \N__40835\
        );

    \I__8789\ : Span4Mux_h
    port map (
            O => \N__40835\,
            I => \N__40832\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__40832\,
            I => buf_data_iac_19
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__40829\,
            I => \n26_adj_1541_cascade_\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__40826\,
            I => \n20837_cascade_\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40820\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40820\,
            I => n22085
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__40817\,
            I => \n22094_cascade_\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40811\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40811\,
            I => \N__40808\
        );

    \I__8780\ : Span12Mux_v
    port map (
            O => \N__40808\,
            I => \N__40805\
        );

    \I__8779\ : Odrv12
    port map (
            O => \N__40805\,
            I => n20828
        );

    \I__8778\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40798\
        );

    \I__8777\ : CascadeMux
    port map (
            O => \N__40801\,
            I => \N__40794\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__40798\,
            I => \N__40789\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40786\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40783\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40780\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40777\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__40789\,
            I => \N__40773\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__40786\,
            I => \N__40770\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40765\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40780\,
            I => \N__40765\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40777\,
            I => \N__40762\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40759\
        );

    \I__8765\ : Span4Mux_v
    port map (
            O => \N__40773\,
            I => \N__40754\
        );

    \I__8764\ : Span4Mux_v
    port map (
            O => \N__40770\,
            I => \N__40751\
        );

    \I__8763\ : Span4Mux_v
    port map (
            O => \N__40765\,
            I => \N__40748\
        );

    \I__8762\ : Span4Mux_v
    port map (
            O => \N__40762\,
            I => \N__40743\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40759\,
            I => \N__40743\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40740\
        );

    \I__8759\ : InMux
    port map (
            O => \N__40757\,
            I => \N__40737\
        );

    \I__8758\ : Span4Mux_h
    port map (
            O => \N__40754\,
            I => \N__40733\
        );

    \I__8757\ : Span4Mux_v
    port map (
            O => \N__40751\,
            I => \N__40730\
        );

    \I__8756\ : Span4Mux_h
    port map (
            O => \N__40748\,
            I => \N__40727\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__40743\,
            I => \N__40724\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40740\,
            I => \N__40721\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40737\,
            I => \N__40718\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40715\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__40733\,
            I => comm_rx_buf_3
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__40730\,
            I => comm_rx_buf_3
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__40727\,
            I => comm_rx_buf_3
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__40724\,
            I => comm_rx_buf_3
        );

    \I__8747\ : Odrv12
    port map (
            O => \N__40721\,
            I => comm_rx_buf_3
        );

    \I__8746\ : Odrv4
    port map (
            O => \N__40718\,
            I => comm_rx_buf_3
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__40715\,
            I => comm_rx_buf_3
        );

    \I__8744\ : CascadeMux
    port map (
            O => \N__40700\,
            I => \n22097_cascade_\
        );

    \I__8743\ : SRMux
    port map (
            O => \N__40697\,
            I => \N__40693\
        );

    \I__8742\ : SRMux
    port map (
            O => \N__40696\,
            I => \N__40690\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__40693\,
            I => \N__40687\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40690\,
            I => \N__40684\
        );

    \I__8739\ : Span4Mux_v
    port map (
            O => \N__40687\,
            I => \N__40681\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__40684\,
            I => \N__40678\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__40681\,
            I => \N__40673\
        );

    \I__8736\ : Span4Mux_h
    port map (
            O => \N__40678\,
            I => \N__40673\
        );

    \I__8735\ : Sp12to4
    port map (
            O => \N__40673\,
            I => \N__40670\
        );

    \I__8734\ : Odrv12
    port map (
            O => \N__40670\,
            I => flagcntwd
        );

    \I__8733\ : CEMux
    port map (
            O => \N__40667\,
            I => \N__40664\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40664\,
            I => n11406
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__40661\,
            I => \N__40658\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40658\,
            I => \N__40655\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__40655\,
            I => \N__40651\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40647\
        );

    \I__8727\ : Span4Mux_v
    port map (
            O => \N__40651\,
            I => \N__40642\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40639\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40647\,
            I => \N__40635\
        );

    \I__8724\ : InMux
    port map (
            O => \N__40646\,
            I => \N__40632\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40645\,
            I => \N__40629\
        );

    \I__8722\ : Span4Mux_h
    port map (
            O => \N__40642\,
            I => \N__40624\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__40639\,
            I => \N__40624\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40638\,
            I => \N__40621\
        );

    \I__8719\ : Span4Mux_v
    port map (
            O => \N__40635\,
            I => \N__40614\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__40632\,
            I => \N__40614\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__40629\,
            I => \N__40611\
        );

    \I__8716\ : Span4Mux_v
    port map (
            O => \N__40624\,
            I => \N__40606\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__40621\,
            I => \N__40606\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40603\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40600\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__40614\,
            I => \N__40596\
        );

    \I__8711\ : Span12Mux_h
    port map (
            O => \N__40611\,
            I => \N__40593\
        );

    \I__8710\ : Span4Mux_v
    port map (
            O => \N__40606\,
            I => \N__40586\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__40603\,
            I => \N__40586\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__40600\,
            I => \N__40586\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40583\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__40596\,
            I => comm_rx_buf_4
        );

    \I__8705\ : Odrv12
    port map (
            O => \N__40593\,
            I => comm_rx_buf_4
        );

    \I__8704\ : Odrv4
    port map (
            O => \N__40586\,
            I => comm_rx_buf_4
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40583\,
            I => comm_rx_buf_4
        );

    \I__8702\ : CascadeMux
    port map (
            O => \N__40574\,
            I => \n30_adj_1539_cascade_\
        );

    \I__8701\ : InMux
    port map (
            O => \N__40571\,
            I => \N__40564\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40564\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__40569\,
            I => \N__40559\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40564\,
            I => \N__40556\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40551\
        );

    \I__8696\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40551\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40548\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__40556\,
            I => \N__40543\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__40551\,
            I => \N__40543\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40538\
        );

    \I__8691\ : Span4Mux_h
    port map (
            O => \N__40543\,
            I => \N__40538\
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__40538\,
            I => comm_cmd_7
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__40535\,
            I => \n20621_cascade_\
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__40532\,
            I => \n25_adj_1619_cascade_\
        );

    \I__8687\ : InMux
    port map (
            O => \N__40529\,
            I => \N__40526\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40526\,
            I => \N__40516\
        );

    \I__8685\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40501\
        );

    \I__8684\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40501\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40501\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40501\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40521\,
            I => \N__40501\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40501\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40501\
        );

    \I__8678\ : Odrv12
    port map (
            O => \N__40516\,
            I => \comm_spi.n16869\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40501\,
            I => \comm_spi.n16869\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40490\
        );

    \I__8674\ : Span4Mux_h
    port map (
            O => \N__40490\,
            I => \N__40487\
        );

    \I__8673\ : Odrv4
    port map (
            O => \N__40487\,
            I => n7_adj_1609
        );

    \I__8672\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40480\
        );

    \I__8671\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40476\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__40480\,
            I => \N__40473\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40470\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40467\
        );

    \I__8667\ : Span12Mux_h
    port map (
            O => \N__40473\,
            I => \N__40464\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40470\,
            I => buf_dds1_11
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__40467\,
            I => buf_dds1_11
        );

    \I__8664\ : Odrv12
    port map (
            O => \N__40464\,
            I => buf_dds1_11
        );

    \I__8663\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40453\
        );

    \I__8662\ : CascadeMux
    port map (
            O => \N__40456\,
            I => \N__40450\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40453\,
            I => \N__40446\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40443\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40449\,
            I => \N__40440\
        );

    \I__8658\ : Span4Mux_v
    port map (
            O => \N__40446\,
            I => \N__40437\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__40443\,
            I => \N__40434\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__40440\,
            I => \N__40427\
        );

    \I__8655\ : Span4Mux_h
    port map (
            O => \N__40437\,
            I => \N__40427\
        );

    \I__8654\ : Span4Mux_v
    port map (
            O => \N__40434\,
            I => \N__40427\
        );

    \I__8653\ : Odrv4
    port map (
            O => \N__40427\,
            I => buf_dds0_11
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__40424\,
            I => \n21506_cascade_\
        );

    \I__8651\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40418\,
            I => \N__40415\
        );

    \I__8649\ : Span12Mux_h
    port map (
            O => \N__40415\,
            I => \N__40412\
        );

    \I__8648\ : Span12Mux_v
    port map (
            O => \N__40412\,
            I => \N__40409\
        );

    \I__8647\ : Odrv12
    port map (
            O => \N__40409\,
            I => n21067
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__40406\,
            I => \N__40403\
        );

    \I__8645\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40400\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40400\,
            I => \N__40397\
        );

    \I__8643\ : Span4Mux_h
    port map (
            O => \N__40397\,
            I => \N__40394\
        );

    \I__8642\ : Span4Mux_v
    port map (
            O => \N__40394\,
            I => \N__40391\
        );

    \I__8641\ : Odrv4
    port map (
            O => \N__40391\,
            I => n23_adj_1538
        );

    \I__8640\ : InMux
    port map (
            O => \N__40388\,
            I => \N__40385\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40385\,
            I => n22028
        );

    \I__8638\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40378\
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__40381\,
            I => \N__40375\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__40378\,
            I => \N__40372\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40375\,
            I => \N__40369\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__40372\,
            I => \N__40366\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40369\,
            I => \N__40363\
        );

    \I__8632\ : Sp12to4
    port map (
            O => \N__40366\,
            I => \N__40359\
        );

    \I__8631\ : Span4Mux_h
    port map (
            O => \N__40363\,
            I => \N__40356\
        );

    \I__8630\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40353\
        );

    \I__8629\ : Span12Mux_h
    port map (
            O => \N__40359\,
            I => \N__40350\
        );

    \I__8628\ : Span4Mux_h
    port map (
            O => \N__40356\,
            I => \N__40347\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__40353\,
            I => buf_adcdata_iac_20
        );

    \I__8626\ : Odrv12
    port map (
            O => \N__40350\,
            I => buf_adcdata_iac_20
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__40347\,
            I => buf_adcdata_iac_20
        );

    \I__8624\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40337\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40334\
        );

    \I__8622\ : Span4Mux_h
    port map (
            O => \N__40334\,
            I => \N__40330\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40333\,
            I => \N__40327\
        );

    \I__8620\ : Span4Mux_v
    port map (
            O => \N__40330\,
            I => \N__40323\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__40327\,
            I => \N__40320\
        );

    \I__8618\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40317\
        );

    \I__8617\ : Span4Mux_v
    port map (
            O => \N__40323\,
            I => \N__40314\
        );

    \I__8616\ : Odrv4
    port map (
            O => \N__40320\,
            I => buf_dds0_12
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40317\,
            I => buf_dds0_12
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__40314\,
            I => buf_dds0_12
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__40307\,
            I => \n22088_cascade_\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40301\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__40301\,
            I => \N__40298\
        );

    \I__8610\ : Span4Mux_h
    port map (
            O => \N__40298\,
            I => \N__40295\
        );

    \I__8609\ : Span4Mux_v
    port map (
            O => \N__40295\,
            I => \N__40290\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40294\,
            I => \N__40287\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40284\
        );

    \I__8606\ : Span4Mux_h
    port map (
            O => \N__40290\,
            I => \N__40281\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40287\,
            I => buf_dds1_12
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__40284\,
            I => buf_dds1_12
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__40281\,
            I => buf_dds1_12
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__40274\,
            I => \n22091_cascade_\
        );

    \I__8601\ : InMux
    port map (
            O => \N__40271\,
            I => \N__40268\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__40268\,
            I => \N__40265\
        );

    \I__8599\ : Span4Mux_v
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8598\ : Sp12to4
    port map (
            O => \N__40262\,
            I => \N__40259\
        );

    \I__8597\ : Odrv12
    port map (
            O => \N__40259\,
            I => n22205
        );

    \I__8596\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40253\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40253\,
            I => n22031
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__40250\,
            I => \n20844_cascade_\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40247\,
            I => \N__40241\
        );

    \I__8592\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40238\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40235\
        );

    \I__8590\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40230\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40241\,
            I => \N__40225\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40225\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40235\,
            I => \N__40222\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40234\,
            I => \N__40219\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40233\,
            I => \N__40216\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__40230\,
            I => \N__40212\
        );

    \I__8583\ : Span4Mux_v
    port map (
            O => \N__40225\,
            I => \N__40205\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__40222\,
            I => \N__40205\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40219\,
            I => \N__40205\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40202\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40215\,
            I => \N__40199\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__40212\,
            I => \N__40188\
        );

    \I__8577\ : Span4Mux_h
    port map (
            O => \N__40205\,
            I => \N__40188\
        );

    \I__8576\ : Span4Mux_v
    port map (
            O => \N__40202\,
            I => \N__40188\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40188\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40185\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40182\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__40188\,
            I => comm_rx_buf_6
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40185\,
            I => comm_rx_buf_6
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__40182\,
            I => comm_rx_buf_6
        );

    \I__8569\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40172\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__40172\,
            I => \N__40167\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40164\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40170\,
            I => \N__40157\
        );

    \I__8565\ : Span4Mux_v
    port map (
            O => \N__40167\,
            I => \N__40152\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40164\,
            I => \N__40152\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40143\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40143\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40143\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40143\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__40157\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__40152\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__40143\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__8556\ : ClkMux
    port map (
            O => \N__40136\,
            I => \N__40128\
        );

    \I__8555\ : ClkMux
    port map (
            O => \N__40135\,
            I => \N__40125\
        );

    \I__8554\ : ClkMux
    port map (
            O => \N__40134\,
            I => \N__40122\
        );

    \I__8553\ : ClkMux
    port map (
            O => \N__40133\,
            I => \N__40113\
        );

    \I__8552\ : ClkMux
    port map (
            O => \N__40132\,
            I => \N__40104\
        );

    \I__8551\ : ClkMux
    port map (
            O => \N__40131\,
            I => \N__40101\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40128\,
            I => \N__40098\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__40125\,
            I => \N__40093\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__40122\,
            I => \N__40093\
        );

    \I__8547\ : ClkMux
    port map (
            O => \N__40121\,
            I => \N__40090\
        );

    \I__8546\ : ClkMux
    port map (
            O => \N__40120\,
            I => \N__40085\
        );

    \I__8545\ : ClkMux
    port map (
            O => \N__40119\,
            I => \N__40082\
        );

    \I__8544\ : ClkMux
    port map (
            O => \N__40118\,
            I => \N__40079\
        );

    \I__8543\ : ClkMux
    port map (
            O => \N__40117\,
            I => \N__40076\
        );

    \I__8542\ : ClkMux
    port map (
            O => \N__40116\,
            I => \N__40073\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__40113\,
            I => \N__40070\
        );

    \I__8540\ : ClkMux
    port map (
            O => \N__40112\,
            I => \N__40067\
        );

    \I__8539\ : ClkMux
    port map (
            O => \N__40111\,
            I => \N__40064\
        );

    \I__8538\ : ClkMux
    port map (
            O => \N__40110\,
            I => \N__40061\
        );

    \I__8537\ : ClkMux
    port map (
            O => \N__40109\,
            I => \N__40057\
        );

    \I__8536\ : ClkMux
    port map (
            O => \N__40108\,
            I => \N__40054\
        );

    \I__8535\ : ClkMux
    port map (
            O => \N__40107\,
            I => \N__40050\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40045\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40042\
        );

    \I__8532\ : Span4Mux_v
    port map (
            O => \N__40098\,
            I => \N__40035\
        );

    \I__8531\ : Span4Mux_h
    port map (
            O => \N__40093\,
            I => \N__40035\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__40090\,
            I => \N__40035\
        );

    \I__8529\ : IoInMux
    port map (
            O => \N__40089\,
            I => \N__40031\
        );

    \I__8528\ : ClkMux
    port map (
            O => \N__40088\,
            I => \N__40028\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__40085\,
            I => \N__40025\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__40082\,
            I => \N__40018\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__40079\,
            I => \N__40018\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__40076\,
            I => \N__40018\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40073\,
            I => \N__40015\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__40070\,
            I => \N__40010\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__40067\,
            I => \N__40010\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__40064\,
            I => \N__40007\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__40061\,
            I => \N__40004\
        );

    \I__8518\ : ClkMux
    port map (
            O => \N__40060\,
            I => \N__40001\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__40057\,
            I => \N__39996\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__40054\,
            I => \N__39996\
        );

    \I__8515\ : ClkMux
    port map (
            O => \N__40053\,
            I => \N__39993\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__39990\
        );

    \I__8513\ : ClkMux
    port map (
            O => \N__40049\,
            I => \N__39987\
        );

    \I__8512\ : ClkMux
    port map (
            O => \N__40048\,
            I => \N__39984\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__40045\,
            I => \N__39981\
        );

    \I__8510\ : Span4Mux_v
    port map (
            O => \N__40042\,
            I => \N__39976\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__40035\,
            I => \N__39976\
        );

    \I__8508\ : ClkMux
    port map (
            O => \N__40034\,
            I => \N__39973\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__40031\,
            I => \N__39970\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__40028\,
            I => \N__39967\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__40025\,
            I => \N__39962\
        );

    \I__8504\ : Span4Mux_v
    port map (
            O => \N__40018\,
            I => \N__39962\
        );

    \I__8503\ : Span4Mux_v
    port map (
            O => \N__40015\,
            I => \N__39957\
        );

    \I__8502\ : Span4Mux_h
    port map (
            O => \N__40010\,
            I => \N__39957\
        );

    \I__8501\ : Span4Mux_v
    port map (
            O => \N__40007\,
            I => \N__39946\
        );

    \I__8500\ : Span4Mux_h
    port map (
            O => \N__40004\,
            I => \N__39946\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__40001\,
            I => \N__39946\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__39996\,
            I => \N__39946\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39993\,
            I => \N__39946\
        );

    \I__8496\ : Span4Mux_v
    port map (
            O => \N__39990\,
            I => \N__39939\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39939\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__39984\,
            I => \N__39939\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__39981\,
            I => \N__39932\
        );

    \I__8492\ : Span4Mux_h
    port map (
            O => \N__39976\,
            I => \N__39932\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39973\,
            I => \N__39932\
        );

    \I__8490\ : Span12Mux_s6_h
    port map (
            O => \N__39970\,
            I => \N__39929\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__39967\,
            I => \N__39926\
        );

    \I__8488\ : Span4Mux_h
    port map (
            O => \N__39962\,
            I => \N__39923\
        );

    \I__8487\ : Span4Mux_v
    port map (
            O => \N__39957\,
            I => \N__39918\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__39946\,
            I => \N__39918\
        );

    \I__8485\ : Span4Mux_v
    port map (
            O => \N__39939\,
            I => \N__39915\
        );

    \I__8484\ : Span4Mux_h
    port map (
            O => \N__39932\,
            I => \N__39912\
        );

    \I__8483\ : Span12Mux_h
    port map (
            O => \N__39929\,
            I => \N__39909\
        );

    \I__8482\ : Span4Mux_h
    port map (
            O => \N__39926\,
            I => \N__39904\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__39923\,
            I => \N__39904\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39899\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__39915\,
            I => \N__39899\
        );

    \I__8478\ : Span4Mux_v
    port map (
            O => \N__39912\,
            I => \N__39896\
        );

    \I__8477\ : Odrv12
    port map (
            O => \N__39909\,
            I => \VDC_CLK\
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__39904\,
            I => \VDC_CLK\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__39899\,
            I => \VDC_CLK\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__39896\,
            I => \VDC_CLK\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39883\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39880\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__39883\,
            I => secclk_cnt_15
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__39880\,
            I => secclk_cnt_15
        );

    \I__8469\ : InMux
    port map (
            O => \N__39875\,
            I => n19523
        );

    \I__8468\ : InMux
    port map (
            O => \N__39872\,
            I => \N__39868\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39871\,
            I => \N__39865\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39868\,
            I => secclk_cnt_16
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39865\,
            I => secclk_cnt_16
        );

    \I__8464\ : InMux
    port map (
            O => \N__39860\,
            I => \bfn_14_20_0_\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39857\,
            I => \N__39853\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39850\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39853\,
            I => secclk_cnt_17
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39850\,
            I => secclk_cnt_17
        );

    \I__8459\ : InMux
    port map (
            O => \N__39845\,
            I => n19525
        );

    \I__8458\ : CascadeMux
    port map (
            O => \N__39842\,
            I => \N__39838\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39835\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39832\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39835\,
            I => secclk_cnt_18
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39832\,
            I => secclk_cnt_18
        );

    \I__8453\ : InMux
    port map (
            O => \N__39827\,
            I => n19526
        );

    \I__8452\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39820\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39817\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__39820\,
            I => secclk_cnt_19
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39817\,
            I => secclk_cnt_19
        );

    \I__8448\ : InMux
    port map (
            O => \N__39812\,
            I => n19527
        );

    \I__8447\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39805\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39802\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39805\,
            I => secclk_cnt_20
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__39802\,
            I => secclk_cnt_20
        );

    \I__8443\ : InMux
    port map (
            O => \N__39797\,
            I => n19528
        );

    \I__8442\ : InMux
    port map (
            O => \N__39794\,
            I => \N__39790\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39787\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39790\,
            I => secclk_cnt_21
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39787\,
            I => secclk_cnt_21
        );

    \I__8438\ : InMux
    port map (
            O => \N__39782\,
            I => n19529
        );

    \I__8437\ : InMux
    port map (
            O => \N__39779\,
            I => n19530
        );

    \I__8436\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39772\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39769\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__39772\,
            I => secclk_cnt_22
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__39769\,
            I => secclk_cnt_22
        );

    \I__8432\ : SRMux
    port map (
            O => \N__39764\,
            I => \N__39760\
        );

    \I__8431\ : SRMux
    port map (
            O => \N__39763\,
            I => \N__39757\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39753\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__39757\,
            I => \N__39750\
        );

    \I__8428\ : SRMux
    port map (
            O => \N__39756\,
            I => \N__39747\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__39753\,
            I => \N__39743\
        );

    \I__8426\ : Span4Mux_h
    port map (
            O => \N__39750\,
            I => \N__39740\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39737\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39746\,
            I => \N__39734\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__39743\,
            I => n14731
        );

    \I__8422\ : Odrv4
    port map (
            O => \N__39740\,
            I => n14731
        );

    \I__8421\ : Odrv4
    port map (
            O => \N__39737\,
            I => n14731
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__39734\,
            I => n14731
        );

    \I__8419\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39721\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39718\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__39721\,
            I => secclk_cnt_7
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39718\,
            I => secclk_cnt_7
        );

    \I__8415\ : InMux
    port map (
            O => \N__39713\,
            I => n19515
        );

    \I__8414\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39706\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39709\,
            I => \N__39703\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39706\,
            I => secclk_cnt_8
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39703\,
            I => secclk_cnt_8
        );

    \I__8410\ : InMux
    port map (
            O => \N__39698\,
            I => \bfn_14_19_0_\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39695\,
            I => \N__39691\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39688\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__39691\,
            I => secclk_cnt_9
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39688\,
            I => secclk_cnt_9
        );

    \I__8405\ : InMux
    port map (
            O => \N__39683\,
            I => n19517
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__39680\,
            I => \N__39676\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39679\,
            I => \N__39673\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39676\,
            I => \N__39670\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__39673\,
            I => secclk_cnt_10
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__39670\,
            I => secclk_cnt_10
        );

    \I__8399\ : InMux
    port map (
            O => \N__39665\,
            I => n19518
        );

    \I__8398\ : InMux
    port map (
            O => \N__39662\,
            I => \N__39658\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39661\,
            I => \N__39655\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__39658\,
            I => secclk_cnt_11
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__39655\,
            I => secclk_cnt_11
        );

    \I__8394\ : InMux
    port map (
            O => \N__39650\,
            I => n19519
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__39647\,
            I => \N__39643\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39640\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39637\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__39640\,
            I => secclk_cnt_12
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__39637\,
            I => secclk_cnt_12
        );

    \I__8388\ : InMux
    port map (
            O => \N__39632\,
            I => n19520
        );

    \I__8387\ : CascadeMux
    port map (
            O => \N__39629\,
            I => \N__39625\
        );

    \I__8386\ : InMux
    port map (
            O => \N__39628\,
            I => \N__39622\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39619\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39622\,
            I => secclk_cnt_13
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__39619\,
            I => secclk_cnt_13
        );

    \I__8382\ : InMux
    port map (
            O => \N__39614\,
            I => n19521
        );

    \I__8381\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39607\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39604\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__39607\,
            I => secclk_cnt_14
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39604\,
            I => secclk_cnt_14
        );

    \I__8377\ : InMux
    port map (
            O => \N__39599\,
            I => n19522
        );

    \I__8376\ : InMux
    port map (
            O => \N__39596\,
            I => n19503
        );

    \I__8375\ : InMux
    port map (
            O => \N__39593\,
            I => n19504
        );

    \I__8374\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39586\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39583\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__39586\,
            I => secclk_cnt_0
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39583\,
            I => secclk_cnt_0
        );

    \I__8370\ : InMux
    port map (
            O => \N__39578\,
            I => \bfn_14_18_0_\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__39575\,
            I => \N__39571\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39568\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39565\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__39568\,
            I => secclk_cnt_1
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__39565\,
            I => secclk_cnt_1
        );

    \I__8364\ : InMux
    port map (
            O => \N__39560\,
            I => n19509
        );

    \I__8363\ : InMux
    port map (
            O => \N__39557\,
            I => \N__39553\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39556\,
            I => \N__39550\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__39553\,
            I => secclk_cnt_2
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39550\,
            I => secclk_cnt_2
        );

    \I__8359\ : InMux
    port map (
            O => \N__39545\,
            I => n19510
        );

    \I__8358\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39538\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39535\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39538\,
            I => secclk_cnt_3
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39535\,
            I => secclk_cnt_3
        );

    \I__8354\ : InMux
    port map (
            O => \N__39530\,
            I => n19511
        );

    \I__8353\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39523\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39520\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39523\,
            I => secclk_cnt_4
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__39520\,
            I => secclk_cnt_4
        );

    \I__8349\ : InMux
    port map (
            O => \N__39515\,
            I => n19512
        );

    \I__8348\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39508\
        );

    \I__8347\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39505\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39508\,
            I => secclk_cnt_5
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__39505\,
            I => secclk_cnt_5
        );

    \I__8344\ : InMux
    port map (
            O => \N__39500\,
            I => n19513
        );

    \I__8343\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39493\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39496\,
            I => \N__39490\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__39493\,
            I => secclk_cnt_6
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__39490\,
            I => secclk_cnt_6
        );

    \I__8339\ : InMux
    port map (
            O => \N__39485\,
            I => n19514
        );

    \I__8338\ : InMux
    port map (
            O => \N__39482\,
            I => \N__39479\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__39479\,
            I => \N__39476\
        );

    \I__8336\ : Odrv12
    port map (
            O => \N__39476\,
            I => n10_adj_1613
        );

    \I__8335\ : InMux
    port map (
            O => \N__39473\,
            I => \bfn_14_17_0_\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39470\,
            I => n19498
        );

    \I__8333\ : InMux
    port map (
            O => \N__39467\,
            I => n19499
        );

    \I__8332\ : InMux
    port map (
            O => \N__39464\,
            I => n19500
        );

    \I__8331\ : InMux
    port map (
            O => \N__39461\,
            I => n19501
        );

    \I__8330\ : InMux
    port map (
            O => \N__39458\,
            I => n19502
        );

    \I__8329\ : InMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__39452\,
            I => n10
        );

    \I__8327\ : CascadeMux
    port map (
            O => \N__39449\,
            I => \N__39446\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39446\,
            I => \N__39443\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__39443\,
            I => \N__39439\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39442\,
            I => \N__39436\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__39439\,
            I => n8_adj_1565
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39436\,
            I => n8_adj_1565
        );

    \I__8321\ : InMux
    port map (
            O => \N__39431\,
            I => \N__39428\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__39428\,
            I => \N__39424\
        );

    \I__8319\ : InMux
    port map (
            O => \N__39427\,
            I => \N__39421\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__39424\,
            I => \N__39418\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39421\,
            I => n7_adj_1564
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__39418\,
            I => n7_adj_1564
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8314\ : CascadeBuf
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__39407\,
            I => \N__39404\
        );

    \I__8312\ : CascadeBuf
    port map (
            O => \N__39404\,
            I => \N__39401\
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__39401\,
            I => \N__39398\
        );

    \I__8310\ : CascadeBuf
    port map (
            O => \N__39398\,
            I => \N__39395\
        );

    \I__8309\ : CascadeMux
    port map (
            O => \N__39395\,
            I => \N__39392\
        );

    \I__8308\ : CascadeBuf
    port map (
            O => \N__39392\,
            I => \N__39389\
        );

    \I__8307\ : CascadeMux
    port map (
            O => \N__39389\,
            I => \N__39386\
        );

    \I__8306\ : CascadeBuf
    port map (
            O => \N__39386\,
            I => \N__39383\
        );

    \I__8305\ : CascadeMux
    port map (
            O => \N__39383\,
            I => \N__39380\
        );

    \I__8304\ : CascadeBuf
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__39377\,
            I => \N__39374\
        );

    \I__8302\ : CascadeBuf
    port map (
            O => \N__39374\,
            I => \N__39371\
        );

    \I__8301\ : CascadeMux
    port map (
            O => \N__39371\,
            I => \N__39368\
        );

    \I__8300\ : CascadeBuf
    port map (
            O => \N__39368\,
            I => \N__39364\
        );

    \I__8299\ : CascadeMux
    port map (
            O => \N__39367\,
            I => \N__39361\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__39364\,
            I => \N__39358\
        );

    \I__8297\ : CascadeBuf
    port map (
            O => \N__39361\,
            I => \N__39355\
        );

    \I__8296\ : CascadeBuf
    port map (
            O => \N__39358\,
            I => \N__39352\
        );

    \I__8295\ : CascadeMux
    port map (
            O => \N__39355\,
            I => \N__39349\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__39352\,
            I => \N__39346\
        );

    \I__8293\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39343\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39346\,
            I => \N__39340\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39337\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__39340\,
            I => \N__39334\
        );

    \I__8289\ : Span12Mux_s10_h
    port map (
            O => \N__39337\,
            I => \N__39331\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__39334\,
            I => \N__39328\
        );

    \I__8287\ : Span12Mux_v
    port map (
            O => \N__39331\,
            I => \N__39325\
        );

    \I__8286\ : Span4Mux_h
    port map (
            O => \N__39328\,
            I => \N__39322\
        );

    \I__8285\ : Odrv12
    port map (
            O => \N__39325\,
            I => \data_index_9_N_216_2\
        );

    \I__8284\ : Odrv4
    port map (
            O => \N__39322\,
            I => \data_index_9_N_216_2\
        );

    \I__8283\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39314\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__39314\,
            I => \N__39310\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39307\
        );

    \I__8280\ : Span4Mux_v
    port map (
            O => \N__39310\,
            I => \N__39304\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39307\,
            I => \N__39301\
        );

    \I__8278\ : Span4Mux_h
    port map (
            O => \N__39304\,
            I => \N__39298\
        );

    \I__8277\ : Span4Mux_v
    port map (
            O => \N__39301\,
            I => \N__39295\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__39298\,
            I => \N__39292\
        );

    \I__8275\ : Span4Mux_h
    port map (
            O => \N__39295\,
            I => \N__39289\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__39292\,
            I => n14_adj_1573
        );

    \I__8273\ : Odrv4
    port map (
            O => \N__39289\,
            I => n14_adj_1573
        );

    \I__8272\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39281\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39281\,
            I => \N__39278\
        );

    \I__8270\ : Span4Mux_h
    port map (
            O => \N__39278\,
            I => \N__39275\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__39275\,
            I => \N__39271\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39268\
        );

    \I__8267\ : Sp12to4
    port map (
            O => \N__39271\,
            I => \N__39263\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__39268\,
            I => \N__39263\
        );

    \I__8265\ : Span12Mux_v
    port map (
            O => \N__39263\,
            I => \N__39260\
        );

    \I__8264\ : Odrv12
    port map (
            O => \N__39260\,
            I => n14_adj_1572
        );

    \I__8263\ : InMux
    port map (
            O => \N__39257\,
            I => \N__39254\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39254\,
            I => \N__39250\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39253\,
            I => \N__39247\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__39250\,
            I => \N__39244\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39247\,
            I => acadc_skipcnt_7
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__39244\,
            I => acadc_skipcnt_7
        );

    \I__8257\ : InMux
    port map (
            O => \N__39239\,
            I => \N__39236\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__39236\,
            I => \N__39232\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39235\,
            I => \N__39229\
        );

    \I__8254\ : Span4Mux_h
    port map (
            O => \N__39232\,
            I => \N__39226\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__39229\,
            I => acadc_skipcnt_2
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__39226\,
            I => acadc_skipcnt_2
        );

    \I__8251\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39218\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__39218\,
            I => n22_adj_1620
        );

    \I__8249\ : CascadeMux
    port map (
            O => \N__39215\,
            I => \N__39212\
        );

    \I__8248\ : InMux
    port map (
            O => \N__39212\,
            I => \N__39209\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__39209\,
            I => \N__39206\
        );

    \I__8246\ : Span4Mux_h
    port map (
            O => \N__39206\,
            I => \N__39203\
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__39203\,
            I => n9_adj_1415
        );

    \I__8244\ : CascadeMux
    port map (
            O => \N__39200\,
            I => \N__39197\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39197\,
            I => \N__39194\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39194\,
            I => \N__39191\
        );

    \I__8241\ : Span4Mux_h
    port map (
            O => \N__39191\,
            I => \N__39187\
        );

    \I__8240\ : InMux
    port map (
            O => \N__39190\,
            I => \N__39184\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__39187\,
            I => \N__39179\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__39184\,
            I => \N__39179\
        );

    \I__8237\ : Span4Mux_v
    port map (
            O => \N__39179\,
            I => \N__39176\
        );

    \I__8236\ : Span4Mux_h
    port map (
            O => \N__39176\,
            I => \N__39173\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__39173\,
            I => n14_adj_1570
        );

    \I__8234\ : InMux
    port map (
            O => \N__39170\,
            I => \N__39167\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__39167\,
            I => \N__39164\
        );

    \I__8232\ : Span12Mux_v
    port map (
            O => \N__39164\,
            I => \N__39161\
        );

    \I__8231\ : Odrv12
    port map (
            O => \N__39161\,
            I => n21048
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__39158\,
            I => \N__39154\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39150\
        );

    \I__8228\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39147\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__39153\,
            I => \N__39144\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__39150\,
            I => \N__39133\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39147\,
            I => \N__39130\
        );

    \I__8224\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39127\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__39143\,
            I => \N__39124\
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__39142\,
            I => \N__39121\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__39141\,
            I => \N__39118\
        );

    \I__8220\ : CascadeMux
    port map (
            O => \N__39140\,
            I => \N__39115\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__39139\,
            I => \N__39112\
        );

    \I__8218\ : CascadeMux
    port map (
            O => \N__39138\,
            I => \N__39109\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__39137\,
            I => \N__39106\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__39136\,
            I => \N__39103\
        );

    \I__8215\ : Span4Mux_h
    port map (
            O => \N__39133\,
            I => \N__39100\
        );

    \I__8214\ : Span4Mux_v
    port map (
            O => \N__39130\,
            I => \N__39097\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__39127\,
            I => \N__39094\
        );

    \I__8212\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39085\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39121\,
            I => \N__39085\
        );

    \I__8210\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39085\
        );

    \I__8209\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39085\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39076\
        );

    \I__8207\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39076\
        );

    \I__8206\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39076\
        );

    \I__8205\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39076\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__39100\,
            I => n10614
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__39097\,
            I => n10614
        );

    \I__8202\ : Odrv12
    port map (
            O => \N__39094\,
            I => n10614
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__39085\,
            I => n10614
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__39076\,
            I => n10614
        );

    \I__8199\ : CEMux
    port map (
            O => \N__39065\,
            I => \N__39062\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__39062\,
            I => \N__39058\
        );

    \I__8197\ : CEMux
    port map (
            O => \N__39061\,
            I => \N__39055\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__39058\,
            I => \N__39052\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__39055\,
            I => \N__39049\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__39052\,
            I => \N__39046\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__39049\,
            I => \N__39043\
        );

    \I__8192\ : Sp12to4
    port map (
            O => \N__39046\,
            I => \N__39040\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__39043\,
            I => n12312
        );

    \I__8190\ : Odrv12
    port map (
            O => \N__39040\,
            I => n12312
        );

    \I__8189\ : IoInMux
    port map (
            O => \N__39035\,
            I => \N__39032\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__39032\,
            I => \N__39029\
        );

    \I__8187\ : IoSpan4Mux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__8186\ : Span4Mux_s2_h
    port map (
            O => \N__39026\,
            I => \N__39023\
        );

    \I__8185\ : Sp12to4
    port map (
            O => \N__39023\,
            I => \N__39020\
        );

    \I__8184\ : Span12Mux_h
    port map (
            O => \N__39020\,
            I => \N__39017\
        );

    \I__8183\ : Span12Mux_v
    port map (
            O => \N__39017\,
            I => \N__39012\
        );

    \I__8182\ : InMux
    port map (
            O => \N__39016\,
            I => \N__39009\
        );

    \I__8181\ : InMux
    port map (
            O => \N__39015\,
            I => \N__39006\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__39012\,
            I => \VDC_RNG0\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__39009\,
            I => \VDC_RNG0\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__39006\,
            I => \VDC_RNG0\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38996\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38996\,
            I => \N__38991\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__38995\,
            I => \N__38988\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38985\
        );

    \I__8173\ : Span4Mux_h
    port map (
            O => \N__38991\,
            I => \N__38982\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38979\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38985\,
            I => \acadc_skipCount_12\
        );

    \I__8170\ : Odrv4
    port map (
            O => \N__38982\,
            I => \acadc_skipCount_12\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__38979\,
            I => \acadc_skipCount_12\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38969\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38969\,
            I => \N__38961\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38958\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38951\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38947\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38944\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38941\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__38961\,
            I => \N__38936\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38936\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38957\,
            I => \N__38925\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38925\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38955\,
            I => \N__38925\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38922\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38951\,
            I => \N__38919\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38916\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38947\,
            I => \N__38913\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__38944\,
            I => \N__38908\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38941\,
            I => \N__38908\
        );

    \I__8150\ : Span4Mux_h
    port map (
            O => \N__38936\,
            I => \N__38905\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38902\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38897\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38897\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38894\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__38925\,
            I => \N__38889\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38889\
        );

    \I__8143\ : Span4Mux_h
    port map (
            O => \N__38919\,
            I => \N__38886\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38916\,
            I => \N__38883\
        );

    \I__8141\ : Span4Mux_h
    port map (
            O => \N__38913\,
            I => \N__38876\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__38908\,
            I => \N__38876\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38905\,
            I => \N__38876\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38902\,
            I => n12383
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38897\,
            I => n12383
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38894\,
            I => n12383
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__38889\,
            I => n12383
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__38886\,
            I => n12383
        );

    \I__8133\ : Odrv12
    port map (
            O => \N__38883\,
            I => n12383
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38876\,
            I => n12383
        );

    \I__8131\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__38858\,
            I => \N__38854\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38851\
        );

    \I__8128\ : Span4Mux_h
    port map (
            O => \N__38854\,
            I => \N__38848\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38851\,
            I => acadc_skipcnt_13
        );

    \I__8126\ : Odrv4
    port map (
            O => \N__38848\,
            I => acadc_skipcnt_13
        );

    \I__8125\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38840\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38840\,
            I => \N__38836\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38832\
        );

    \I__8122\ : Span4Mux_v
    port map (
            O => \N__38836\,
            I => \N__38829\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38826\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38832\,
            I => \acadc_skipCount_13\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__38829\,
            I => \acadc_skipCount_13\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38826\,
            I => \acadc_skipCount_13\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38819\,
            I => \N__38816\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38816\,
            I => n14
        );

    \I__8115\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38810\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38810\,
            I => \N__38806\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38803\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__38806\,
            I => \N__38800\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38803\,
            I => acadc_skipcnt_1
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__38800\,
            I => acadc_skipcnt_1
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__38795\,
            I => \N__38792\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38789\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38789\,
            I => \N__38785\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38782\
        );

    \I__8105\ : Span4Mux_v
    port map (
            O => \N__38785\,
            I => \N__38779\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__38782\,
            I => acadc_skipcnt_4
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__38779\,
            I => acadc_skipcnt_4
        );

    \I__8102\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38771\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__38771\,
            I => n18_adj_1611
        );

    \I__8100\ : InMux
    port map (
            O => \N__38768\,
            I => \N__38764\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38767\,
            I => \N__38761\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38764\,
            I => \N__38756\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__38761\,
            I => \N__38756\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__38756\,
            I => \N__38752\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38749\
        );

    \I__8094\ : Span4Mux_h
    port map (
            O => \N__38752\,
            I => \N__38746\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38749\,
            I => data_index_4
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__38746\,
            I => data_index_4
        );

    \I__8091\ : InMux
    port map (
            O => \N__38741\,
            I => \N__38735\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38740\,
            I => \N__38735\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__38735\,
            I => \N__38732\
        );

    \I__8088\ : Span4Mux_v
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__38729\,
            I => n7_adj_1560
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__38726\,
            I => \N__38722\
        );

    \I__8085\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38717\
        );

    \I__8084\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38717\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__38717\,
            I => n8_adj_1561
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__8081\ : CascadeBuf
    port map (
            O => \N__38711\,
            I => \N__38708\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__8079\ : CascadeBuf
    port map (
            O => \N__38705\,
            I => \N__38702\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__38702\,
            I => \N__38699\
        );

    \I__8077\ : CascadeBuf
    port map (
            O => \N__38699\,
            I => \N__38696\
        );

    \I__8076\ : CascadeMux
    port map (
            O => \N__38696\,
            I => \N__38693\
        );

    \I__8075\ : CascadeBuf
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__38690\,
            I => \N__38687\
        );

    \I__8073\ : CascadeBuf
    port map (
            O => \N__38687\,
            I => \N__38684\
        );

    \I__8072\ : CascadeMux
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__8071\ : CascadeBuf
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__8069\ : CascadeBuf
    port map (
            O => \N__38675\,
            I => \N__38672\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__38672\,
            I => \N__38669\
        );

    \I__8067\ : CascadeBuf
    port map (
            O => \N__38669\,
            I => \N__38665\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__38668\,
            I => \N__38662\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__38665\,
            I => \N__38659\
        );

    \I__8064\ : CascadeBuf
    port map (
            O => \N__38662\,
            I => \N__38656\
        );

    \I__8063\ : CascadeBuf
    port map (
            O => \N__38659\,
            I => \N__38653\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__38656\,
            I => \N__38650\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__38653\,
            I => \N__38647\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38644\
        );

    \I__8059\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38641\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__38644\,
            I => \N__38638\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__38641\,
            I => \N__38635\
        );

    \I__8056\ : Span12Mux_s11_h
    port map (
            O => \N__38638\,
            I => \N__38632\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__38635\,
            I => \N__38629\
        );

    \I__8054\ : Span12Mux_v
    port map (
            O => \N__38632\,
            I => \N__38626\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__38629\,
            I => \N__38623\
        );

    \I__8052\ : Odrv12
    port map (
            O => \N__38626\,
            I => \data_index_9_N_216_4\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__38623\,
            I => \data_index_9_N_216_4\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__38615\,
            I => n22013
        );

    \I__8048\ : CascadeMux
    port map (
            O => \N__38612\,
            I => \n12441_cascade_\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__38609\,
            I => \n8_adj_1567_cascade_\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38602\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38605\,
            I => \N__38599\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38602\,
            I => \N__38594\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38599\,
            I => \N__38594\
        );

    \I__8042\ : Span4Mux_v
    port map (
            O => \N__38594\,
            I => \N__38590\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38587\
        );

    \I__8040\ : Span4Mux_h
    port map (
            O => \N__38590\,
            I => \N__38584\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__38587\,
            I => data_index_1
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__38584\,
            I => data_index_1
        );

    \I__8037\ : CascadeMux
    port map (
            O => \N__38579\,
            I => \N__38575\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38568\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38564\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38552\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38549\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38572\,
            I => \N__38544\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38544\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__38568\,
            I => \N__38541\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38538\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__38564\,
            I => \N__38535\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38532\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38529\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38561\,
            I => \N__38524\
        );

    \I__8024\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38524\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38521\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38516\
        );

    \I__8021\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38516\
        );

    \I__8020\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38511\
        );

    \I__8019\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38511\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__38552\,
            I => \N__38502\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38549\,
            I => \N__38502\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38502\
        );

    \I__8015\ : Span4Mux_h
    port map (
            O => \N__38541\,
            I => \N__38502\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__38538\,
            I => \N__38497\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__38535\,
            I => \N__38497\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__38532\,
            I => n11835
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38529\,
            I => n11835
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38524\,
            I => n11835
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__38521\,
            I => n11835
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__38516\,
            I => n11835
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__38511\,
            I => n11835
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__38502\,
            I => n11835
        );

    \I__8005\ : Odrv4
    port map (
            O => \N__38497\,
            I => n11835
        );

    \I__8004\ : InMux
    port map (
            O => \N__38480\,
            I => \N__38476\
        );

    \I__8003\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38476\,
            I => \N__38467\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38464\
        );

    \I__8000\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38461\
        );

    \I__7999\ : InMux
    port map (
            O => \N__38471\,
            I => \N__38456\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38456\
        );

    \I__7997\ : Span4Mux_h
    port map (
            O => \N__38467\,
            I => \N__38445\
        );

    \I__7996\ : Span4Mux_h
    port map (
            O => \N__38464\,
            I => \N__38440\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38461\,
            I => \N__38440\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38456\,
            I => \N__38437\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38434\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38431\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38426\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38426\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38423\
        );

    \I__7988\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38416\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38416\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38416\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__38445\,
            I => n16763
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__38440\,
            I => n16763
        );

    \I__7983\ : Odrv12
    port map (
            O => \N__38437\,
            I => n16763
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__38434\,
            I => n16763
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38431\,
            I => n16763
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38426\,
            I => n16763
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__38423\,
            I => n16763
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38416\,
            I => n16763
        );

    \I__7977\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38395\
        );

    \I__7976\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38389\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38385\
        );

    \I__7973\ : Span4Mux_h
    port map (
            O => \N__38389\,
            I => \N__38382\
        );

    \I__7972\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38379\
        );

    \I__7971\ : Span12Mux_h
    port map (
            O => \N__38385\,
            I => \N__38376\
        );

    \I__7970\ : Span4Mux_h
    port map (
            O => \N__38382\,
            I => \N__38373\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__38379\,
            I => buf_dds1_1
        );

    \I__7968\ : Odrv12
    port map (
            O => \N__38376\,
            I => buf_dds1_1
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__38373\,
            I => buf_dds1_1
        );

    \I__7966\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__38363\,
            I => \N__38360\
        );

    \I__7964\ : Span4Mux_h
    port map (
            O => \N__38360\,
            I => \N__38356\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38353\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__38356\,
            I => \N__38347\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38344\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__38347\,
            I => \N__38341\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__38344\,
            I => buf_adcdata_iac_14
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__38341\,
            I => buf_adcdata_iac_14
        );

    \I__7956\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38333\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__38333\,
            I => \N__38330\
        );

    \I__7954\ : Span4Mux_h
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__38327\,
            I => n16
        );

    \I__7952\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__7950\ : Odrv12
    port map (
            O => \N__38318\,
            I => n20953
        );

    \I__7949\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38312\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__38312\,
            I => \N__38308\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38305\
        );

    \I__7946\ : Odrv12
    port map (
            O => \N__38308\,
            I => \buf_readRTD_3\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__38305\,
            I => \buf_readRTD_3\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__38297\,
            I => n20879
        );

    \I__7942\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__38291\,
            I => \N__38287\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__38290\,
            I => \N__38283\
        );

    \I__7939\ : Span4Mux_h
    port map (
            O => \N__38287\,
            I => \N__38280\
        );

    \I__7938\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38277\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38283\,
            I => \N__38274\
        );

    \I__7936\ : Span4Mux_h
    port map (
            O => \N__38280\,
            I => \N__38271\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38277\,
            I => \N__38268\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38274\,
            I => \N__38263\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__38271\,
            I => \N__38263\
        );

    \I__7932\ : Odrv4
    port map (
            O => \N__38268\,
            I => buf_adcdata_vac_11
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__38263\,
            I => buf_adcdata_vac_11
        );

    \I__7930\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38255\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38255\,
            I => \N__38252\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__38252\,
            I => \N__38249\
        );

    \I__7927\ : Span4Mux_h
    port map (
            O => \N__38249\,
            I => \N__38245\
        );

    \I__7926\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38242\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__38245\,
            I => buf_adcdata_vdc_11
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38242\,
            I => buf_adcdata_vdc_11
        );

    \I__7923\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38234\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__38234\,
            I => n19_adj_1513
        );

    \I__7921\ : CascadeMux
    port map (
            O => \N__38231\,
            I => \n22178_cascade_\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__38228\,
            I => \n22181_cascade_\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__38225\,
            I => \n30_adj_1511_cascade_\
        );

    \I__7918\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__38219\,
            I => \N__38215\
        );

    \I__7916\ : CascadeMux
    port map (
            O => \N__38218\,
            I => \N__38212\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__38215\,
            I => \N__38209\
        );

    \I__7914\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38206\
        );

    \I__7913\ : Sp12to4
    port map (
            O => \N__38209\,
            I => \N__38203\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__38206\,
            I => data_idxvec_4
        );

    \I__7911\ : Odrv12
    port map (
            O => \N__38203\,
            I => data_idxvec_4
        );

    \I__7910\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38195\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__38195\,
            I => n26_adj_1510
        );

    \I__7908\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38189\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__38189\,
            I => n19_adj_1509
        );

    \I__7906\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38183\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__38183\,
            I => \N__38179\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__38182\,
            I => \N__38176\
        );

    \I__7903\ : Sp12to4
    port map (
            O => \N__38179\,
            I => \N__38173\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38170\
        );

    \I__7901\ : Odrv12
    port map (
            O => \N__38173\,
            I => \buf_readRTD_4\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38170\,
            I => \buf_readRTD_4\
        );

    \I__7899\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38162\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__38162\,
            I => \N__38158\
        );

    \I__7897\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38155\
        );

    \I__7896\ : Span4Mux_h
    port map (
            O => \N__38158\,
            I => \N__38152\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__38155\,
            I => \N__38149\
        );

    \I__7894\ : Span4Mux_h
    port map (
            O => \N__38152\,
            I => \N__38145\
        );

    \I__7893\ : Span4Mux_v
    port map (
            O => \N__38149\,
            I => \N__38142\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38139\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__38145\,
            I => \N__38136\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__38142\,
            I => \N__38133\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38139\,
            I => buf_adcdata_iac_12
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__38136\,
            I => buf_adcdata_iac_12
        );

    \I__7887\ : Odrv4
    port map (
            O => \N__38133\,
            I => buf_adcdata_iac_12
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__38126\,
            I => \n22010_cascade_\
        );

    \I__7885\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38120\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__38120\,
            I => \N__38117\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__38117\,
            I => \N__38114\
        );

    \I__7882\ : Span4Mux_h
    port map (
            O => \N__38114\,
            I => \N__38111\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__38111\,
            I => n16_adj_1508
        );

    \I__7880\ : InMux
    port map (
            O => \N__38108\,
            I => \N__38105\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__38105\,
            I => \N__38102\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__38102\,
            I => \N__38098\
        );

    \I__7877\ : CascadeMux
    port map (
            O => \N__38101\,
            I => \N__38095\
        );

    \I__7876\ : Span4Mux_h
    port map (
            O => \N__38098\,
            I => \N__38092\
        );

    \I__7875\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38089\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__38092\,
            I => buf_adcdata_vdc_14
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__38089\,
            I => buf_adcdata_vdc_14
        );

    \I__7872\ : InMux
    port map (
            O => \N__38084\,
            I => \N__38081\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__38081\,
            I => \N__38078\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__38078\,
            I => \N__38073\
        );

    \I__7869\ : CascadeMux
    port map (
            O => \N__38077\,
            I => \N__38070\
        );

    \I__7868\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38067\
        );

    \I__7867\ : Span4Mux_v
    port map (
            O => \N__38073\,
            I => \N__38064\
        );

    \I__7866\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38061\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__38067\,
            I => \N__38056\
        );

    \I__7864\ : Span4Mux_h
    port map (
            O => \N__38064\,
            I => \N__38056\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__38061\,
            I => buf_adcdata_vac_14
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__38056\,
            I => buf_adcdata_vac_14
        );

    \I__7861\ : InMux
    port map (
            O => \N__38051\,
            I => \N__38048\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__38048\,
            I => \N__38045\
        );

    \I__7859\ : Span12Mux_h
    port map (
            O => \N__38045\,
            I => \N__38041\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38038\
        );

    \I__7857\ : Odrv12
    port map (
            O => \N__38041\,
            I => \buf_readRTD_6\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__38038\,
            I => \buf_readRTD_6\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__38033\,
            I => \n19_cascade_\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38027\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__38027\,
            I => \N__38024\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__38024\,
            I => n20954
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__7850\ : InMux
    port map (
            O => \N__38018\,
            I => \N__38015\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__38015\,
            I => \N__38010\
        );

    \I__7848\ : InMux
    port map (
            O => \N__38014\,
            I => \N__38007\
        );

    \I__7847\ : InMux
    port map (
            O => \N__38013\,
            I => \N__38004\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__38010\,
            I => \N__38001\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__38007\,
            I => \N__37998\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__38004\,
            I => \acadc_skipCount_6\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__38001\,
            I => \acadc_skipCount_6\
        );

    \I__7842\ : Odrv12
    port map (
            O => \N__37998\,
            I => \acadc_skipCount_6\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37991\,
            I => \N__37988\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__37988\,
            I => n20929
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__37985\,
            I => \N__37982\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37978\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37975\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37978\,
            I => \N__37972\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37975\,
            I => \N__37966\
        );

    \I__7834\ : Span4Mux_h
    port map (
            O => \N__37972\,
            I => \N__37963\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37958\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37970\,
            I => \N__37958\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37955\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__37966\,
            I => \N__37952\
        );

    \I__7829\ : Span4Mux_h
    port map (
            O => \N__37963\,
            I => \N__37947\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37958\,
            I => \N__37947\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__37955\,
            I => \N__37944\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__37952\,
            I => \N__37941\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__37947\,
            I => \N__37938\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__37944\,
            I => comm_buf_1_3
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__37941\,
            I => comm_buf_1_3
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__37938\,
            I => comm_buf_1_3
        );

    \I__7821\ : InMux
    port map (
            O => \N__37931\,
            I => \N__37926\
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__37930\,
            I => \N__37923\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__37929\,
            I => \N__37920\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37917\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37912\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37912\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__37917\,
            I => \acadc_skipCount_3\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37912\,
            I => \acadc_skipCount_3\
        );

    \I__7813\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \n20884_cascade_\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37901\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__37901\,
            I => \N__37898\
        );

    \I__7810\ : Span4Mux_h
    port map (
            O => \N__37898\,
            I => \N__37895\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__37895\,
            I => \N__37892\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37892\,
            I => n20878
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__37889\,
            I => \n22124_cascade_\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37883\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37883\,
            I => n22127
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__37880\,
            I => \N__37877\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37873\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37870\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37873\,
            I => \N__37865\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37865\
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__37865\,
            I => data_idxvec_3
        );

    \I__7798\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37859\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37859\,
            I => \N__37856\
        );

    \I__7796\ : Span4Mux_v
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7795\ : Span4Mux_h
    port map (
            O => \N__37853\,
            I => \N__37850\
        );

    \I__7794\ : Span4Mux_h
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__7793\ : Span4Mux_h
    port map (
            O => \N__37847\,
            I => \N__37844\
        );

    \I__7792\ : Odrv4
    port map (
            O => \N__37844\,
            I => buf_data_iac_11
        );

    \I__7791\ : CascadeMux
    port map (
            O => \N__37841\,
            I => \n26_adj_1514_cascade_\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37835\,
            I => n20885
        );

    \I__7788\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37829\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__37829\,
            I => \N__37826\
        );

    \I__7786\ : Odrv12
    port map (
            O => \N__37826\,
            I => comm_buf_3_3
        );

    \I__7785\ : InMux
    port map (
            O => \N__37823\,
            I => \N__37820\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37820\,
            I => \N__37817\
        );

    \I__7783\ : Span4Mux_h
    port map (
            O => \N__37817\,
            I => \N__37814\
        );

    \I__7782\ : Sp12to4
    port map (
            O => \N__37814\,
            I => \N__37811\
        );

    \I__7781\ : Odrv12
    port map (
            O => \N__37811\,
            I => comm_buf_2_3
        );

    \I__7780\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37805\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37805\,
            I => n2_adj_1590
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__37802\,
            I => \n21102_cascade_\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37799\,
            I => \N__37796\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__37796\,
            I => n21_adj_1618
        );

    \I__7775\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37790\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37790\,
            I => n16_adj_1599
        );

    \I__7773\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37783\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__37786\,
            I => \N__37780\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37783\,
            I => \N__37777\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37774\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__37777\,
            I => \N__37771\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__37774\,
            I => data_idxvec_6
        );

    \I__7767\ : Odrv4
    port map (
            O => \N__37771\,
            I => data_idxvec_6
        );

    \I__7766\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37763\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37760\
        );

    \I__7764\ : Span4Mux_h
    port map (
            O => \N__37760\,
            I => \N__37757\
        );

    \I__7763\ : Span4Mux_h
    port map (
            O => \N__37757\,
            I => \N__37754\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__37754\,
            I => buf_data_iac_14
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__37751\,
            I => \n26_adj_1505_cascade_\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__37748\,
            I => \n20930_cascade_\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__37745\,
            I => \n21962_cascade_\
        );

    \I__7758\ : CascadeMux
    port map (
            O => \N__37742\,
            I => \n21965_cascade_\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37736\,
            I => \N__37733\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__37733\,
            I => \N__37730\
        );

    \I__7754\ : Span4Mux_v
    port map (
            O => \N__37730\,
            I => \N__37727\
        );

    \I__7753\ : Span4Mux_v
    port map (
            O => \N__37727\,
            I => \N__37724\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__37724\,
            I => buf_data_vac_12
        );

    \I__7751\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37718\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37718\,
            I => \N__37715\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__37715\,
            I => \N__37712\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__37712\,
            I => comm_buf_4_4
        );

    \I__7747\ : InMux
    port map (
            O => \N__37709\,
            I => \N__37706\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37706\,
            I => \N__37703\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__37703\,
            I => \N__37700\
        );

    \I__7744\ : Span4Mux_v
    port map (
            O => \N__37700\,
            I => \N__37697\
        );

    \I__7743\ : Span4Mux_h
    port map (
            O => \N__37697\,
            I => \N__37694\
        );

    \I__7742\ : Span4Mux_h
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__7741\ : Odrv4
    port map (
            O => \N__37691\,
            I => buf_data_vac_11
        );

    \I__7740\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37685\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__7738\ : Span4Mux_h
    port map (
            O => \N__37682\,
            I => \N__37679\
        );

    \I__7737\ : Span4Mux_h
    port map (
            O => \N__37679\,
            I => \N__37676\
        );

    \I__7736\ : Span4Mux_v
    port map (
            O => \N__37676\,
            I => \N__37673\
        );

    \I__7735\ : Span4Mux_v
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__7734\ : Odrv4
    port map (
            O => \N__37670\,
            I => buf_data_vac_10
        );

    \I__7733\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37664\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37661\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__7730\ : Span4Mux_h
    port map (
            O => \N__37658\,
            I => \N__37655\
        );

    \I__7729\ : Span4Mux_v
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__7728\ : Span4Mux_v
    port map (
            O => \N__37652\,
            I => \N__37649\
        );

    \I__7727\ : Odrv4
    port map (
            O => \N__37649\,
            I => buf_data_vac_9
        );

    \I__7726\ : CEMux
    port map (
            O => \N__37646\,
            I => \N__37643\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37643\,
            I => \N__37640\
        );

    \I__7724\ : Span4Mux_h
    port map (
            O => \N__37640\,
            I => \N__37637\
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__37637\,
            I => n12194
        );

    \I__7722\ : SRMux
    port map (
            O => \N__37634\,
            I => \N__37631\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__37631\,
            I => \N__37628\
        );

    \I__7720\ : Span4Mux_h
    port map (
            O => \N__37628\,
            I => \N__37625\
        );

    \I__7719\ : Odrv4
    port map (
            O => \N__37625\,
            I => n14794
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__37622\,
            I => \n1_adj_1589_cascade_\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37615\
        );

    \I__7716\ : InMux
    port map (
            O => \N__37618\,
            I => \N__37612\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__37615\,
            I => \N__37609\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37612\,
            I => comm_buf_6_3
        );

    \I__7713\ : Odrv4
    port map (
            O => \N__37609\,
            I => comm_buf_6_3
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__37604\,
            I => \n21296_cascade_\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37598\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__37598\,
            I => n22154
        );

    \I__7709\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37592\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37592\,
            I => comm_buf_4_3
        );

    \I__7707\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37586\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__37586\,
            I => \N__37583\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__37583\,
            I => \N__37580\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__37580\,
            I => comm_buf_5_3
        );

    \I__7703\ : InMux
    port map (
            O => \N__37577\,
            I => \N__37574\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__37574\,
            I => n4_adj_1591
        );

    \I__7701\ : CascadeMux
    port map (
            O => \N__37571\,
            I => \N__37568\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37565\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37565\,
            I => comm_buf_2_0
        );

    \I__7698\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37559\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37556\
        );

    \I__7696\ : Odrv12
    port map (
            O => \N__37556\,
            I => comm_buf_3_0
        );

    \I__7695\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37550\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37550\,
            I => n2
        );

    \I__7693\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37544\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7691\ : Span4Mux_v
    port map (
            O => \N__37541\,
            I => \N__37538\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__37538\,
            I => comm_buf_5_0
        );

    \I__7689\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37532\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__37532\,
            I => n20970
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__37529\,
            I => \n4_adj_1507_cascade_\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__37523\,
            I => n21980
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__37520\,
            I => \n21116_cascade_\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37513\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37509\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37513\,
            I => \N__37506\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37503\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37509\,
            I => \N__37500\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__37506\,
            I => \N__37495\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37495\
        );

    \I__7676\ : Span12Mux_h
    port map (
            O => \N__37500\,
            I => \N__37492\
        );

    \I__7675\ : Span4Mux_v
    port map (
            O => \N__37495\,
            I => \N__37489\
        );

    \I__7674\ : Span12Mux_v
    port map (
            O => \N__37492\,
            I => \N__37486\
        );

    \I__7673\ : Span4Mux_v
    port map (
            O => \N__37489\,
            I => \N__37483\
        );

    \I__7672\ : Odrv12
    port map (
            O => \N__37486\,
            I => n10713
        );

    \I__7671\ : Odrv4
    port map (
            O => \N__37483\,
            I => n10713
        );

    \I__7670\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__37475\,
            I => n12_adj_1602
        );

    \I__7668\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__7666\ : Span12Mux_h
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7665\ : Span12Mux_v
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__7664\ : Odrv12
    port map (
            O => \N__37460\,
            I => buf_data_vac_8
        );

    \I__7663\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__37454\,
            I => comm_buf_4_0
        );

    \I__7661\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37448\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37445\
        );

    \I__7659\ : Span4Mux_h
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7657\ : Span4Mux_v
    port map (
            O => \N__37439\,
            I => \N__37436\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__37436\,
            I => buf_data_vac_15
        );

    \I__7655\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37430\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37427\
        );

    \I__7653\ : Span12Mux_h
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7652\ : Odrv12
    port map (
            O => \N__37424\,
            I => buf_data_vac_14
        );

    \I__7651\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__37418\,
            I => \N__37415\
        );

    \I__7649\ : Span4Mux_h
    port map (
            O => \N__37415\,
            I => \N__37412\
        );

    \I__7648\ : Span4Mux_v
    port map (
            O => \N__37412\,
            I => \N__37409\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__37406\,
            I => buf_data_vac_13
        );

    \I__7645\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37400\,
            I => \N__37397\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__37397\,
            I => \N__37394\
        );

    \I__7642\ : Span4Mux_h
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__37388\,
            I => buf_data_vac_23
        );

    \I__7639\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7637\ : Span4Mux_v
    port map (
            O => \N__37379\,
            I => \N__37376\
        );

    \I__7636\ : Span4Mux_h
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7635\ : Odrv4
    port map (
            O => \N__37373\,
            I => buf_data_vac_22
        );

    \I__7634\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37367\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__37364\,
            I => \N__37361\
        );

    \I__7631\ : Span4Mux_h
    port map (
            O => \N__37361\,
            I => \N__37358\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__37358\,
            I => buf_data_vac_21
        );

    \I__7629\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__37352\,
            I => \N__37349\
        );

    \I__7627\ : Span4Mux_h
    port map (
            O => \N__37349\,
            I => \N__37346\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__37343\,
            I => buf_data_vac_19
        );

    \I__7624\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37334\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7621\ : Span4Mux_v
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7619\ : Odrv4
    port map (
            O => \N__37325\,
            I => buf_data_vac_18
        );

    \I__7618\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37319\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37316\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__37316\,
            I => \N__37313\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__37313\,
            I => \N__37310\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__37307\,
            I => buf_data_vac_17
        );

    \I__7612\ : CEMux
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37298\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__37298\,
            I => \N__37295\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__37295\,
            I => n12152
        );

    \I__7608\ : SRMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__37289\,
            I => n14787
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__37286\,
            I => \n1_cascade_\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__37283\,
            I => \n30_adj_1535_cascade_\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__37280\,
            I => \N__37277\
        );

    \I__7603\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37273\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37270\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__37273\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__37270\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__7599\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37261\
        );

    \I__7598\ : InMux
    port map (
            O => \N__37264\,
            I => \N__37258\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37261\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__37258\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__37253\,
            I => \N__37249\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__37252\,
            I => \N__37246\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37243\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37240\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37237\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37240\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__37237\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__7588\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37228\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37225\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__37228\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__37225\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__37220\,
            I => \ADC_VDC.genclk.n21211_cascade_\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__37217\,
            I => \N__37213\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37210\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37207\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N__37202\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37207\,
            I => \N__37202\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__37202\,
            I => \ADC_VDC.genclk.n21205\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37195\
        );

    \I__7576\ : InMux
    port map (
            O => \N__37198\,
            I => \N__37192\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__37195\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__37192\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37183\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37180\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37183\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37180\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__37175\,
            I => \N__37171\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37168\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37165\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__37168\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__37165\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__7564\ : CascadeMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37153\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37150\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__37153\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37150\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__7559\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__37142\,
            I => \ADC_VDC.genclk.n26_adj_1408\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__7556\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37132\
        );

    \I__7555\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37129\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__37132\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__37129\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37120\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37117\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37120\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__37117\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__37112\,
            I => \N__37108\
        );

    \I__7547\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37105\
        );

    \I__7546\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37102\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__37105\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__37102\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__7543\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37093\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37090\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__37093\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37090\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__7539\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__37082\,
            I => \ADC_VDC.genclk.n28_adj_1407\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__7536\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37072\
        );

    \I__7535\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37069\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__37072\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__37069\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37057\
        );

    \I__7530\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37054\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__37057\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__37054\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__37049\,
            I => \N__37045\
        );

    \I__7526\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37042\
        );

    \I__7525\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37039\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__37042\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__37039\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7521\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37027\
        );

    \I__7520\ : InMux
    port map (
            O => \N__37030\,
            I => \N__37024\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__37027\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__37024\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__7517\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__37016\,
            I => \ADC_VDC.genclk.n27_adj_1409\
        );

    \I__7515\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__7513\ : Span12Mux_h
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7512\ : Odrv12
    port map (
            O => \N__37004\,
            I => buf_data_vac_16
        );

    \I__7511\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7509\ : Span4Mux_v
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7508\ : Span4Mux_h
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__36989\,
            I => buf_data_vac_20
        );

    \I__7506\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7504\ : Odrv12
    port map (
            O => \N__36980\,
            I => comm_buf_3_4
        );

    \I__7503\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36974\,
            I => n28_adj_1621
        );

    \I__7501\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36968\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36968\,
            I => n14_adj_1592
        );

    \I__7499\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36961\
        );

    \I__7498\ : CascadeMux
    port map (
            O => \N__36964\,
            I => \N__36958\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36961\,
            I => \N__36955\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36951\
        );

    \I__7495\ : Span4Mux_v
    port map (
            O => \N__36955\,
            I => \N__36948\
        );

    \I__7494\ : CascadeMux
    port map (
            O => \N__36954\,
            I => \N__36945\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36951\,
            I => \N__36942\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__36948\,
            I => \N__36939\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36936\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__36942\,
            I => \N__36931\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__36939\,
            I => \N__36931\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36936\,
            I => buf_dds1_14
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__36931\,
            I => buf_dds1_14
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__36926\,
            I => \N__36922\
        );

    \I__7485\ : CascadeMux
    port map (
            O => \N__36925\,
            I => \N__36919\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36922\,
            I => \N__36916\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36913\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__36916\,
            I => \N__36910\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36906\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36910\,
            I => \N__36903\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36900\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__36906\,
            I => \N__36897\
        );

    \I__7477\ : Span4Mux_v
    port map (
            O => \N__36903\,
            I => \N__36894\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36900\,
            I => buf_dds0_14
        );

    \I__7475\ : Odrv4
    port map (
            O => \N__36897\,
            I => buf_dds0_14
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36894\,
            I => buf_dds0_14
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__36887\,
            I => \n22115_cascade_\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36884\,
            I => \N__36881\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36878\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__36878\,
            I => \N__36875\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__36872\,
            I => n22163
        );

    \I__7467\ : IoInMux
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36866\,
            I => \N__36862\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36859\
        );

    \I__7464\ : Span4Mux_s0_h
    port map (
            O => \N__36862\,
            I => \N__36856\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36859\,
            I => \N__36853\
        );

    \I__7462\ : Sp12to4
    port map (
            O => \N__36856\,
            I => \N__36850\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__36853\,
            I => \N__36847\
        );

    \I__7460\ : Span12Mux_v
    port map (
            O => \N__36850\,
            I => \N__36844\
        );

    \I__7459\ : Span4Mux_v
    port map (
            O => \N__36847\,
            I => \N__36840\
        );

    \I__7458\ : Span12Mux_h
    port map (
            O => \N__36844\,
            I => \N__36837\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36834\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__36840\,
            I => \N__36831\
        );

    \I__7455\ : Odrv12
    port map (
            O => \N__36837\,
            I => \VAC_FLT0\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36834\,
            I => \VAC_FLT0\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__36831\,
            I => \VAC_FLT0\
        );

    \I__7452\ : CascadeMux
    port map (
            O => \N__36824\,
            I => \N__36821\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36817\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36814\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36817\,
            I => \N__36811\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36808\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__36811\,
            I => \N__36805\
        );

    \I__7446\ : Span4Mux_v
    port map (
            O => \N__36808\,
            I => \N__36802\
        );

    \I__7445\ : Span4Mux_v
    port map (
            O => \N__36805\,
            I => \N__36799\
        );

    \I__7444\ : Span4Mux_v
    port map (
            O => \N__36802\,
            I => \N__36796\
        );

    \I__7443\ : Sp12to4
    port map (
            O => \N__36799\,
            I => \N__36790\
        );

    \I__7442\ : Sp12to4
    port map (
            O => \N__36796\,
            I => \N__36790\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36787\
        );

    \I__7440\ : Span12Mux_h
    port map (
            O => \N__36790\,
            I => \N__36784\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36787\,
            I => buf_adcdata_iac_22
        );

    \I__7438\ : Odrv12
    port map (
            O => \N__36784\,
            I => buf_adcdata_iac_22
        );

    \I__7437\ : InMux
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36776\,
            I => n22112
        );

    \I__7435\ : CascadeMux
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__36755\,
            I => n21037
        );

    \I__7428\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36749\,
            I => \N__36746\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7425\ : Span4Mux_v
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__36740\,
            I => n23_adj_1534
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__36737\,
            I => \n22070_cascade_\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__36731\,
            I => n20856
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__36728\,
            I => \n22073_cascade_\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__36725\,
            I => \N__36721\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36710\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36710\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36702\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36702\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36693\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36693\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36693\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36693\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36710\,
            I => \N__36690\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36687\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36680\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36680\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36702\,
            I => \N__36677\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36669\
        );

    \I__7404\ : Span4Mux_v
    port map (
            O => \N__36690\,
            I => \N__36669\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__36687\,
            I => \N__36666\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36686\,
            I => \N__36661\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36685\,
            I => \N__36661\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36680\,
            I => \N__36658\
        );

    \I__7399\ : Span4Mux_v
    port map (
            O => \N__36677\,
            I => \N__36655\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36648\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36648\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36648\
        );

    \I__7395\ : Odrv4
    port map (
            O => \N__36669\,
            I => \eis_end_N_725\
        );

    \I__7394\ : Odrv12
    port map (
            O => \N__36666\,
            I => \eis_end_N_725\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__36661\,
            I => \eis_end_N_725\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__36658\,
            I => \eis_end_N_725\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__36655\,
            I => \eis_end_N_725\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36648\,
            I => \eis_end_N_725\
        );

    \I__7389\ : CEMux
    port map (
            O => \N__36635\,
            I => \N__36631\
        );

    \I__7388\ : CEMux
    port map (
            O => \N__36634\,
            I => \N__36628\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__36631\,
            I => \N__36624\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__36628\,
            I => \N__36621\
        );

    \I__7385\ : CEMux
    port map (
            O => \N__36627\,
            I => \N__36618\
        );

    \I__7384\ : Span4Mux_v
    port map (
            O => \N__36624\,
            I => \N__36614\
        );

    \I__7383\ : Span4Mux_h
    port map (
            O => \N__36621\,
            I => \N__36609\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36609\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36606\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__36614\,
            I => n11670
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__36609\,
            I => n11670
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36606\,
            I => n11670
        );

    \I__7377\ : SRMux
    port map (
            O => \N__36599\,
            I => \N__36595\
        );

    \I__7376\ : SRMux
    port map (
            O => \N__36598\,
            I => \N__36592\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36595\,
            I => n14687
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__36592\,
            I => n14687
        );

    \I__7373\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36583\
        );

    \I__7372\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36579\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36576\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36582\,
            I => \N__36573\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__36579\,
            I => \N__36569\
        );

    \I__7368\ : Span4Mux_v
    port map (
            O => \N__36576\,
            I => \N__36564\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__36573\,
            I => \N__36564\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36572\,
            I => \N__36561\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__36569\,
            I => \N__36558\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__36564\,
            I => \N__36555\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__36561\,
            I => n10733
        );

    \I__7362\ : Odrv4
    port map (
            O => \N__36558\,
            I => n10733
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__36555\,
            I => n10733
        );

    \I__7360\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36544\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36540\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__36544\,
            I => \N__36537\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36534\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__36540\,
            I => \N__36531\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__36537\,
            I => buf_dds0_5
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__36534\,
            I => buf_dds0_5
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__36531\,
            I => buf_dds0_5
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__36524\,
            I => \n27_adj_1551_cascade_\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36518\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36518\,
            I => n25
        );

    \I__7349\ : CascadeMux
    port map (
            O => \N__36515\,
            I => \n19608_cascade_\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36509\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__36509\,
            I => n10_adj_1594
        );

    \I__7346\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36503\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__36503\,
            I => n26_adj_1543
        );

    \I__7344\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36497\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36493\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36496\,
            I => \N__36490\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__36493\,
            I => \N__36487\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36490\,
            I => acadc_skipcnt_15
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__36487\,
            I => acadc_skipcnt_15
        );

    \I__7338\ : InMux
    port map (
            O => \N__36482\,
            I => \N__36478\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36481\,
            I => \N__36475\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__36478\,
            I => \N__36472\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__36475\,
            I => acadc_skipcnt_9
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__36472\,
            I => acadc_skipcnt_9
        );

    \I__7333\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36464\,
            I => n21
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__36461\,
            I => \n24_adj_1537_cascade_\
        );

    \I__7330\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36455\,
            I => n23_adj_1624
        );

    \I__7328\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36449\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__36449\,
            I => n30
        );

    \I__7326\ : SRMux
    port map (
            O => \N__36446\,
            I => \N__36443\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36443\,
            I => \N__36440\
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__36440\,
            I => n20789
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36428\
        );

    \I__7321\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36425\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36422\
        );

    \I__7319\ : CascadeMux
    port map (
            O => \N__36431\,
            I => \N__36411\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36428\,
            I => \N__36408\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36425\,
            I => \N__36405\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__36422\,
            I => \N__36402\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36399\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36420\,
            I => \N__36396\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36391\
        );

    \I__7312\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36391\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36382\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36382\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36382\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36382\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36379\
        );

    \I__7306\ : Span4Mux_v
    port map (
            O => \N__36408\,
            I => \N__36370\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__36405\,
            I => \N__36370\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__36402\,
            I => \N__36370\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__36399\,
            I => \N__36370\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36396\,
            I => eis_state_0
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__36391\,
            I => eis_state_0
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36382\,
            I => eis_state_0
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__36379\,
            I => eis_state_0
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__36370\,
            I => eis_state_0
        );

    \I__7297\ : InMux
    port map (
            O => \N__36359\,
            I => \N__36356\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__36353\,
            I => \N__36349\
        );

    \I__7294\ : SRMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__36349\,
            I => \N__36339\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36346\,
            I => \N__36339\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36330\
        );

    \I__7290\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36330\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__36339\,
            I => \N__36327\
        );

    \I__7288\ : SRMux
    port map (
            O => \N__36338\,
            I => \N__36324\
        );

    \I__7287\ : InMux
    port map (
            O => \N__36337\,
            I => \N__36321\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36316\
        );

    \I__7285\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36316\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36330\,
            I => \N__36313\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__36327\,
            I => acadc_rst
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__36324\,
            I => acadc_rst
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__36321\,
            I => acadc_rst
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36316\,
            I => acadc_rst
        );

    \I__7279\ : Odrv12
    port map (
            O => \N__36313\,
            I => acadc_rst
        );

    \I__7278\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36299\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36296\
        );

    \I__7276\ : Sp12to4
    port map (
            O => \N__36296\,
            I => \N__36292\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36288\
        );

    \I__7274\ : Span12Mux_v
    port map (
            O => \N__36292\,
            I => \N__36285\
        );

    \I__7273\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36282\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__36288\,
            I => buf_dds1_5
        );

    \I__7271\ : Odrv12
    port map (
            O => \N__36285\,
            I => buf_dds1_5
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__36282\,
            I => buf_dds1_5
        );

    \I__7269\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36271\
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__36274\,
            I => \N__36268\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36271\,
            I => \N__36265\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36262\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__36265\,
            I => \N__36259\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__36262\,
            I => data_idxvec_14
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__36259\,
            I => data_idxvec_14
        );

    \I__7262\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36250\
        );

    \I__7261\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__36247\,
            I => acadc_skipcnt_5
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__36244\,
            I => acadc_skipcnt_5
        );

    \I__7257\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36236\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__36236\,
            I => \N__36232\
        );

    \I__7255\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36229\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__36232\,
            I => \N__36226\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__36229\,
            I => acadc_skipcnt_3
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__36226\,
            I => acadc_skipcnt_3
        );

    \I__7251\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36218\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__36218\,
            I => \N__36214\
        );

    \I__7249\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36211\
        );

    \I__7248\ : Span4Mux_h
    port map (
            O => \N__36214\,
            I => \N__36208\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36211\,
            I => acadc_skipcnt_8
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__36208\,
            I => acadc_skipcnt_8
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__36203\,
            I => \n20_adj_1617_cascade_\
        );

    \I__7244\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36197\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__36197\,
            I => n17_adj_1612
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__36194\,
            I => \n26_adj_1640_cascade_\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36185\
        );

    \I__7240\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36185\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__36185\,
            I => n31
        );

    \I__7238\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36177\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36174\
        );

    \I__7236\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36171\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36166\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__36174\,
            I => \N__36166\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36171\,
            I => \N__36161\
        );

    \I__7232\ : Span4Mux_v
    port map (
            O => \N__36166\,
            I => \N__36161\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__36161\,
            I => data_index_2
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__36158\,
            I => \n11_cascade_\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__36155\,
            I => \n21099_cascade_\
        );

    \I__7228\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__36149\,
            I => n13
        );

    \I__7226\ : CEMux
    port map (
            O => \N__36146\,
            I => \N__36143\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__36143\,
            I => \N__36139\
        );

    \I__7224\ : CEMux
    port map (
            O => \N__36142\,
            I => \N__36136\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__36139\,
            I => \N__36131\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__36136\,
            I => \N__36131\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__36131\,
            I => n11760
        );

    \I__7220\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36125\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__36125\,
            I => n17430
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__36122\,
            I => \N__36115\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__36121\,
            I => \N__36112\
        );

    \I__7216\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36106\
        );

    \I__7215\ : InMux
    port map (
            O => \N__36119\,
            I => \N__36106\
        );

    \I__7214\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36103\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36096\
        );

    \I__7212\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36096\
        );

    \I__7211\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36096\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__36106\,
            I => \N__36093\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__36103\,
            I => acadc_dtrig_v
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36096\,
            I => acadc_dtrig_v
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__36093\,
            I => acadc_dtrig_v
        );

    \I__7206\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36072\
        );

    \I__7205\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36072\
        );

    \I__7204\ : InMux
    port map (
            O => \N__36084\,
            I => \N__36072\
        );

    \I__7203\ : InMux
    port map (
            O => \N__36083\,
            I => \N__36072\
        );

    \I__7202\ : InMux
    port map (
            O => \N__36082\,
            I => \N__36067\
        );

    \I__7201\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36067\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__36072\,
            I => acadc_dtrig_i
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__36067\,
            I => acadc_dtrig_i
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__7197\ : InMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__36056\,
            I => \N__36053\
        );

    \I__7195\ : Span4Mux_v
    port map (
            O => \N__36053\,
            I => \N__36050\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__36050\,
            I => n4_adj_1569
        );

    \I__7193\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36043\
        );

    \I__7192\ : InMux
    port map (
            O => \N__36046\,
            I => \N__36040\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__36043\,
            I => \N__36034\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__36040\,
            I => \N__36034\
        );

    \I__7189\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36031\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__36031\,
            I => data_index_3
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__36028\,
            I => data_index_3
        );

    \I__7185\ : InMux
    port map (
            O => \N__36023\,
            I => \N__36020\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__36020\,
            I => n8_adj_1563
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__36017\,
            I => \n8_adj_1563_cascade_\
        );

    \I__7182\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36008\
        );

    \I__7181\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36008\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__36005\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__36005\,
            I => n7_adj_1562
        );

    \I__7178\ : CascadeMux
    port map (
            O => \N__36002\,
            I => \N__35999\
        );

    \I__7177\ : CascadeBuf
    port map (
            O => \N__35999\,
            I => \N__35996\
        );

    \I__7176\ : CascadeMux
    port map (
            O => \N__35996\,
            I => \N__35993\
        );

    \I__7175\ : CascadeBuf
    port map (
            O => \N__35993\,
            I => \N__35990\
        );

    \I__7174\ : CascadeMux
    port map (
            O => \N__35990\,
            I => \N__35987\
        );

    \I__7173\ : CascadeBuf
    port map (
            O => \N__35987\,
            I => \N__35984\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__35984\,
            I => \N__35981\
        );

    \I__7171\ : CascadeBuf
    port map (
            O => \N__35981\,
            I => \N__35978\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__35978\,
            I => \N__35975\
        );

    \I__7169\ : CascadeBuf
    port map (
            O => \N__35975\,
            I => \N__35972\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__35972\,
            I => \N__35969\
        );

    \I__7167\ : CascadeBuf
    port map (
            O => \N__35969\,
            I => \N__35966\
        );

    \I__7166\ : CascadeMux
    port map (
            O => \N__35966\,
            I => \N__35963\
        );

    \I__7165\ : CascadeBuf
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7164\ : CascadeMux
    port map (
            O => \N__35960\,
            I => \N__35956\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__35959\,
            I => \N__35953\
        );

    \I__7162\ : CascadeBuf
    port map (
            O => \N__35956\,
            I => \N__35950\
        );

    \I__7161\ : CascadeBuf
    port map (
            O => \N__35953\,
            I => \N__35947\
        );

    \I__7160\ : CascadeMux
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__35947\,
            I => \N__35941\
        );

    \I__7158\ : CascadeBuf
    port map (
            O => \N__35944\,
            I => \N__35938\
        );

    \I__7157\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35935\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__35938\,
            I => \N__35932\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35935\,
            I => \N__35929\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35926\
        );

    \I__7153\ : Span4Mux_v
    port map (
            O => \N__35929\,
            I => \N__35923\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35926\,
            I => \N__35920\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__35923\,
            I => \N__35917\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__35917\,
            I => \N__35911\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__35914\,
            I => \N__35908\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__35911\,
            I => \N__35905\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__35908\,
            I => \N__35902\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__35905\,
            I => \data_index_9_N_216_3\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35902\,
            I => \data_index_9_N_216_3\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__35888\,
            I => n16598
        );

    \I__7139\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35882\,
            I => \N__35879\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35879\,
            I => n20957
        );

    \I__7136\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35873\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__35873\,
            I => \N__35870\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__35870\,
            I => \N__35864\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35869\,
            I => \N__35861\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__35868\,
            I => \N__35852\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__35867\,
            I => \N__35848\
        );

    \I__7130\ : Span4Mux_h
    port map (
            O => \N__35864\,
            I => \N__35844\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35861\,
            I => \N__35841\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35836\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35836\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35831\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35831\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35828\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35817\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35817\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35817\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35817\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35817\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__35844\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__35841\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35836\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__35831\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35828\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35817\,
            I => \DTRIG_N_919_adj_1451\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35800\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35803\,
            I => \N__35796\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35793\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35781\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35776\
        );

    \I__7107\ : Span12Mux_h
    port map (
            O => \N__35793\,
            I => \N__35776\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35769\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35769\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35769\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35766\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35761\
        );

    \I__7101\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35761\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35754\
        );

    \I__7099\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35754\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35754\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35781\,
            I => adc_state_1_adj_1417
        );

    \I__7096\ : Odrv12
    port map (
            O => \N__35776\,
            I => adc_state_1_adj_1417
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35769\,
            I => adc_state_1_adj_1417
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35766\,
            I => adc_state_1_adj_1417
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35761\,
            I => adc_state_1_adj_1417
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35754\,
            I => adc_state_1_adj_1417
        );

    \I__7091\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35738\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35735\
        );

    \I__7089\ : Span4Mux_v
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__7088\ : Sp12to4
    port map (
            O => \N__35732\,
            I => \N__35729\
        );

    \I__7087\ : Span12Mux_h
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__7086\ : Span12Mux_v
    port map (
            O => \N__35726\,
            I => \N__35723\
        );

    \I__7085\ : Odrv12
    port map (
            O => \N__35723\,
            I => \ICE_GPMO_0\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35713\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35710\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__35713\,
            I => \N__35707\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35710\,
            I => \N__35704\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__35707\,
            I => \N__35699\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__35704\,
            I => \N__35699\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__35699\,
            I => \N__35694\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35691\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35688\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__35694\,
            I => auxmode
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35691\,
            I => auxmode
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__35688\,
            I => auxmode
        );

    \I__7071\ : CascadeMux
    port map (
            O => \N__35681\,
            I => \acadc_rst_cascade_\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35670\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35665\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35673\,
            I => \N__35665\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__35670\,
            I => tacadc_rst
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35665\,
            I => tacadc_rst
        );

    \I__7064\ : InMux
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35654\
        );

    \I__7062\ : Span4Mux_h
    port map (
            O => \N__35654\,
            I => \N__35650\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35647\
        );

    \I__7060\ : Odrv4
    port map (
            O => \N__35650\,
            I => \buf_readRTD_7\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__35647\,
            I => \buf_readRTD_7\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35639\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__35639\,
            I => \N__35636\
        );

    \I__7056\ : Span4Mux_v
    port map (
            O => \N__35636\,
            I => \N__35633\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__35633\,
            I => n19_adj_1502
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__35630\,
            I => \n24_adj_1622_cascade_\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35624\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__35624\,
            I => \N__35621\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__35621\,
            I => \N__35618\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__35618\,
            I => \N__35615\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__35615\,
            I => \N__35611\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35614\,
            I => \N__35608\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__35611\,
            I => buf_adcdata_vdc_12
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__35608\,
            I => buf_adcdata_vdc_12
        );

    \I__7045\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35600\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__35600\,
            I => \N__35597\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__35597\,
            I => \N__35594\
        );

    \I__7042\ : Span4Mux_h
    port map (
            O => \N__35594\,
            I => \N__35590\
        );

    \I__7041\ : InMux
    port map (
            O => \N__35593\,
            I => \N__35586\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__35590\,
            I => \N__35583\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35580\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__35586\,
            I => buf_adcdata_vac_12
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__35583\,
            I => buf_adcdata_vac_12
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__35580\,
            I => buf_adcdata_vac_12
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \n35_cascade_\
        );

    \I__7034\ : SRMux
    port map (
            O => \N__35570\,
            I => \N__35563\
        );

    \I__7033\ : SRMux
    port map (
            O => \N__35569\,
            I => \N__35559\
        );

    \I__7032\ : SRMux
    port map (
            O => \N__35568\,
            I => \N__35555\
        );

    \I__7031\ : SRMux
    port map (
            O => \N__35567\,
            I => \N__35551\
        );

    \I__7030\ : SRMux
    port map (
            O => \N__35566\,
            I => \N__35547\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35543\
        );

    \I__7028\ : SRMux
    port map (
            O => \N__35562\,
            I => \N__35540\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35536\
        );

    \I__7026\ : SRMux
    port map (
            O => \N__35558\,
            I => \N__35533\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35555\,
            I => \N__35530\
        );

    \I__7024\ : SRMux
    port map (
            O => \N__35554\,
            I => \N__35527\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35524\
        );

    \I__7022\ : SRMux
    port map (
            O => \N__35550\,
            I => \N__35521\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35518\
        );

    \I__7020\ : SRMux
    port map (
            O => \N__35546\,
            I => \N__35515\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__35543\,
            I => \N__35510\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35510\
        );

    \I__7017\ : SRMux
    port map (
            O => \N__35539\,
            I => \N__35507\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__35536\,
            I => \N__35501\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35533\,
            I => \N__35501\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__35530\,
            I => \N__35498\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35527\,
            I => \N__35495\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__35524\,
            I => \N__35492\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35489\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__35518\,
            I => \N__35484\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__35515\,
            I => \N__35484\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__35510\,
            I => \N__35479\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__35507\,
            I => \N__35479\
        );

    \I__7006\ : SRMux
    port map (
            O => \N__35506\,
            I => \N__35476\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__35501\,
            I => \N__35473\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__35498\,
            I => \N__35468\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__35495\,
            I => \N__35468\
        );

    \I__7002\ : Span4Mux_v
    port map (
            O => \N__35492\,
            I => \N__35463\
        );

    \I__7001\ : Span4Mux_h
    port map (
            O => \N__35489\,
            I => \N__35463\
        );

    \I__7000\ : Span4Mux_v
    port map (
            O => \N__35484\,
            I => \N__35458\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35458\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35455\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__35473\,
            I => \N__35452\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__35468\,
            I => \N__35443\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__35463\,
            I => \N__35443\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__35458\,
            I => \N__35443\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__35455\,
            I => \N__35443\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__35452\,
            I => \N__35440\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__35443\,
            I => \N__35437\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__35440\,
            I => \iac_raw_buf_N_735\
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__35437\,
            I => \iac_raw_buf_N_735\
        );

    \I__6988\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__35426\,
            I => n17_adj_1645
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__35423\,
            I => \N__35413\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__35422\,
            I => \N__35397\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35387\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35382\
        );

    \I__6981\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35382\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35377\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35377\
        );

    \I__6978\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35373\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35358\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35412\,
            I => \N__35353\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35353\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35348\
        );

    \I__6973\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35348\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35332\
        );

    \I__6971\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35332\
        );

    \I__6970\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35332\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35332\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35404\,
            I => \N__35321\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35321\
        );

    \I__6966\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35321\
        );

    \I__6965\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35321\
        );

    \I__6964\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35321\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35397\,
            I => \N__35316\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35307\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35307\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35307\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35307\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35298\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35298\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35390\,
            I => \N__35298\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35291\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35382\,
            I => \N__35291\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35291\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35288\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__35373\,
            I => \N__35285\
        );

    \I__6950\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35270\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35270\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35270\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35270\
        );

    \I__6946\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35270\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35367\,
            I => \N__35270\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35270\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35259\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35259\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35259\
        );

    \I__6940\ : InMux
    port map (
            O => \N__35362\,
            I => \N__35259\
        );

    \I__6939\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35259\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35256\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35253\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__35348\,
            I => \N__35250\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35243\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35346\,
            I => \N__35243\
        );

    \I__6933\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35243\
        );

    \I__6932\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35234\
        );

    \I__6931\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35234\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35234\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35234\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35229\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35229\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35320\,
            I => \N__35224\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35224\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35316\,
            I => \N__35219\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__35307\,
            I => \N__35219\
        );

    \I__6922\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35211\
        );

    \I__6921\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35208\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__35298\,
            I => \N__35205\
        );

    \I__6919\ : Span4Mux_v
    port map (
            O => \N__35291\,
            I => \N__35202\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35197\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__35285\,
            I => \N__35197\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35192\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35192\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__35256\,
            I => \N__35185\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__35253\,
            I => \N__35185\
        );

    \I__6912\ : Span4Mux_v
    port map (
            O => \N__35250\,
            I => \N__35185\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__35243\,
            I => \N__35178\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35178\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__35229\,
            I => \N__35178\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__35224\,
            I => \N__35175\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__35219\,
            I => \N__35172\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35158\
        );

    \I__6905\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35158\
        );

    \I__6904\ : InMux
    port map (
            O => \N__35216\,
            I => \N__35158\
        );

    \I__6903\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35153\
        );

    \I__6902\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35153\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35150\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__35208\,
            I => \N__35147\
        );

    \I__6899\ : Span4Mux_h
    port map (
            O => \N__35205\,
            I => \N__35140\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__35202\,
            I => \N__35140\
        );

    \I__6897\ : Span4Mux_h
    port map (
            O => \N__35197\,
            I => \N__35140\
        );

    \I__6896\ : Span4Mux_v
    port map (
            O => \N__35192\,
            I => \N__35134\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__35185\,
            I => \N__35134\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__35178\,
            I => \N__35131\
        );

    \I__6893\ : Span4Mux_h
    port map (
            O => \N__35175\,
            I => \N__35125\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__35172\,
            I => \N__35122\
        );

    \I__6891\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35115\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35115\
        );

    \I__6889\ : InMux
    port map (
            O => \N__35169\,
            I => \N__35115\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35112\
        );

    \I__6887\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35109\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35106\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35103\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__35158\,
            I => \N__35096\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35153\,
            I => \N__35096\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__35150\,
            I => \N__35096\
        );

    \I__6881\ : Span12Mux_v
    port map (
            O => \N__35147\,
            I => \N__35091\
        );

    \I__6880\ : Sp12to4
    port map (
            O => \N__35140\,
            I => \N__35091\
        );

    \I__6879\ : InMux
    port map (
            O => \N__35139\,
            I => \N__35088\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__35134\,
            I => \N__35083\
        );

    \I__6877\ : Span4Mux_h
    port map (
            O => \N__35131\,
            I => \N__35083\
        );

    \I__6876\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35076\
        );

    \I__6875\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35076\
        );

    \I__6874\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35076\
        );

    \I__6873\ : Span4Mux_v
    port map (
            O => \N__35125\,
            I => \N__35069\
        );

    \I__6872\ : Span4Mux_h
    port map (
            O => \N__35122\,
            I => \N__35069\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35115\,
            I => \N__35069\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__35112\,
            I => adc_state_0
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__35109\,
            I => adc_state_0
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__35106\,
            I => adc_state_0
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__35103\,
            I => adc_state_0
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__35096\,
            I => adc_state_0
        );

    \I__6865\ : Odrv12
    port map (
            O => \N__35091\,
            I => adc_state_0
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35088\,
            I => adc_state_0
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__35083\,
            I => adc_state_0
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35076\,
            I => adc_state_0
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__35069\,
            I => adc_state_0
        );

    \I__6860\ : InMux
    port map (
            O => \N__35048\,
            I => \N__35045\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35045\,
            I => \N__35041\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35038\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__35041\,
            I => \N__35035\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__35032\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__35035\,
            I => \N__35026\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__35032\,
            I => \N__35021\
        );

    \I__6853\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35014\
        );

    \I__6852\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35009\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35009\
        );

    \I__6850\ : Span4Mux_h
    port map (
            O => \N__35026\,
            I => \N__35005\
        );

    \I__6849\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35000\
        );

    \I__6848\ : InMux
    port map (
            O => \N__35024\,
            I => \N__35000\
        );

    \I__6847\ : Span4Mux_h
    port map (
            O => \N__35021\,
            I => \N__34997\
        );

    \I__6846\ : InMux
    port map (
            O => \N__35020\,
            I => \N__34988\
        );

    \I__6845\ : InMux
    port map (
            O => \N__35019\,
            I => \N__34988\
        );

    \I__6844\ : InMux
    port map (
            O => \N__35018\,
            I => \N__34988\
        );

    \I__6843\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34988\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34983\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__34983\
        );

    \I__6840\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34980\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__35005\,
            I => adc_state_1
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__35000\,
            I => adc_state_1
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__34997\,
            I => adc_state_1
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34988\,
            I => adc_state_1
        );

    \I__6835\ : Odrv12
    port map (
            O => \N__34983\,
            I => adc_state_1
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34980\,
            I => adc_state_1
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__34967\,
            I => \N__34964\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34961\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34956\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34953\
        );

    \I__6829\ : CascadeMux
    port map (
            O => \N__34959\,
            I => \N__34950\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__34956\,
            I => \N__34946\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__34953\,
            I => \N__34942\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34933\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34949\,
            I => \N__34933\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__34946\,
            I => \N__34930\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__34945\,
            I => \N__34927\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__34942\,
            I => \N__34921\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34918\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34913\
        );

    \I__6819\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34913\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34910\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34933\,
            I => \N__34905\
        );

    \I__6816\ : Span4Mux_h
    port map (
            O => \N__34930\,
            I => \N__34905\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34927\,
            I => \N__34896\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34896\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34896\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34896\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__34921\,
            I => \N__34893\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34888\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34888\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34910\,
            I => \DTRIG_N_919\
        );

    \I__6807\ : Odrv4
    port map (
            O => \N__34905\,
            I => \DTRIG_N_919\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34896\,
            I => \DTRIG_N_919\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__34893\,
            I => \DTRIG_N_919\
        );

    \I__6804\ : Odrv12
    port map (
            O => \N__34888\,
            I => \DTRIG_N_919\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__34877\,
            I => \N__34874\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34871\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__6800\ : Odrv12
    port map (
            O => \N__34868\,
            I => n8
        );

    \I__6799\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34861\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__34864\,
            I => \N__34858\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34855\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34852\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__34855\,
            I => \N__34849\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34852\,
            I => \N__34846\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__34849\,
            I => n11354
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__34846\,
            I => n11354
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \n10534_cascade_\
        );

    \I__6790\ : CascadeMux
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34831\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__34834\,
            I => \N__34826\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34823\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34820\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34815\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34815\
        );

    \I__6783\ : Span4Mux_h
    port map (
            O => \N__34823\,
            I => \N__34812\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34809\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34815\,
            I => \N__34806\
        );

    \I__6780\ : Span4Mux_h
    port map (
            O => \N__34812\,
            I => \N__34803\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__34809\,
            I => n20670
        );

    \I__6778\ : Odrv12
    port map (
            O => \N__34806\,
            I => n20670
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__34803\,
            I => n20670
        );

    \I__6776\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34792\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__34792\,
            I => \N__34786\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34789\,
            I => \N__34783\
        );

    \I__6772\ : Span12Mux_h
    port map (
            O => \N__34786\,
            I => \N__34780\
        );

    \I__6771\ : Span12Mux_v
    port map (
            O => \N__34783\,
            I => \N__34777\
        );

    \I__6770\ : Odrv12
    port map (
            O => \N__34780\,
            I => n20672
        );

    \I__6769\ : Odrv12
    port map (
            O => \N__34777\,
            I => n20672
        );

    \I__6768\ : CascadeMux
    port map (
            O => \N__34772\,
            I => \N__34769\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34762\
        );

    \I__6765\ : CascadeMux
    port map (
            O => \N__34765\,
            I => \N__34758\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__34762\,
            I => \N__34755\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34750\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34750\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__34755\,
            I => cmd_rdadctmp_9
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34750\,
            I => cmd_rdadctmp_9
        );

    \I__6759\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34742\,
            I => \N__34738\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34735\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__34738\,
            I => \N__34731\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__34735\,
            I => \N__34728\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34725\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__34731\,
            I => \N__34720\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__34728\,
            I => \N__34720\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34725\,
            I => buf_adcdata_vac_1
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__34720\,
            I => buf_adcdata_vac_1
        );

    \I__6749\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__6747\ : Odrv4
    port map (
            O => \N__34709\,
            I => n20840
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__34706\,
            I => \N__34703\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34698\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34693\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34693\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__34698\,
            I => cmd_rdadctmp_21
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34693\,
            I => cmd_rdadctmp_21
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__34688\,
            I => \N__34683\
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__34687\,
            I => \N__34680\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__34686\,
            I => \N__34677\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34674\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34671\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34668\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__34674\,
            I => cmd_rdadctmp_20
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__34671\,
            I => cmd_rdadctmp_20
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__34668\,
            I => cmd_rdadctmp_20
        );

    \I__6731\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34641\
        );

    \I__6730\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34641\
        );

    \I__6729\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34641\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34638\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34631\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34631\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34631\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34628\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34625\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34618\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34609\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34609\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34609\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34609\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34606\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__34638\,
            I => \N__34599\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__34631\,
            I => \N__34599\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34599\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34625\,
            I => \N__34596\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34588\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34588\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34585\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34580\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34577\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__34609\,
            I => \N__34574\
        );

    \I__6706\ : Span4Mux_v
    port map (
            O => \N__34606\,
            I => \N__34569\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__34599\,
            I => \N__34569\
        );

    \I__6704\ : Span4Mux_v
    port map (
            O => \N__34596\,
            I => \N__34566\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34563\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34558\
        );

    \I__6701\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34558\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34588\,
            I => \N__34553\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34553\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34548\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34583\,
            I => \N__34548\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__34580\,
            I => \N__34543\
        );

    \I__6695\ : Span12Mux_s9_v
    port map (
            O => \N__34577\,
            I => \N__34543\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__34574\,
            I => \N__34538\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__34569\,
            I => \N__34538\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__34566\,
            I => \N__34535\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__34563\,
            I => n20590
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__34558\,
            I => n20590
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__34553\,
            I => n20590
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__34548\,
            I => n20590
        );

    \I__6687\ : Odrv12
    port map (
            O => \N__34543\,
            I => n20590
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__34538\,
            I => n20590
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__34535\,
            I => n20590
        );

    \I__6684\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34515\
        );

    \I__6683\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34512\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__34518\,
            I => \N__34509\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34506\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34512\,
            I => \N__34503\
        );

    \I__6679\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34500\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34497\
        );

    \I__6677\ : Span4Mux_v
    port map (
            O => \N__34503\,
            I => \N__34494\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__34500\,
            I => cmd_rdadctmp_19
        );

    \I__6675\ : Odrv4
    port map (
            O => \N__34497\,
            I => cmd_rdadctmp_19
        );

    \I__6674\ : Odrv4
    port map (
            O => \N__34494\,
            I => cmd_rdadctmp_19
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__34487\,
            I => \N__34484\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34479\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34476\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__34482\,
            I => \N__34473\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__34479\,
            I => \N__34468\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34468\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34465\
        );

    \I__6666\ : Odrv12
    port map (
            O => \N__34468\,
            I => cmd_rdadctmp_25
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__34465\,
            I => cmd_rdadctmp_25
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__34460\,
            I => \N__34457\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34447\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34447\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34444\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34441\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34436\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34433\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34419\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34444\,
            I => \N__34419\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34416\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34411\
        );

    \I__6653\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34411\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34405\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34405\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34402\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34399\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34396\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34393\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34388\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34388\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34383\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34383\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34377\
        );

    \I__6641\ : Span4Mux_h
    port map (
            O => \N__34419\,
            I => \N__34370\
        );

    \I__6640\ : Span4Mux_v
    port map (
            O => \N__34416\,
            I => \N__34370\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34411\,
            I => \N__34370\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34367\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__34405\,
            I => \N__34362\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34402\,
            I => \N__34362\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__34399\,
            I => \N__34357\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34357\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__34393\,
            I => \N__34350\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__34388\,
            I => \N__34350\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__34383\,
            I => \N__34350\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34343\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34343\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34380\,
            I => \N__34343\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34340\
        );

    \I__6626\ : Span4Mux_v
    port map (
            O => \N__34370\,
            I => \N__34329\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34367\,
            I => \N__34326\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__34362\,
            I => \N__34317\
        );

    \I__6623\ : Span4Mux_v
    port map (
            O => \N__34357\,
            I => \N__34317\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__34350\,
            I => \N__34317\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34343\,
            I => \N__34317\
        );

    \I__6620\ : Span4Mux_v
    port map (
            O => \N__34340\,
            I => \N__34314\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34305\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34305\
        );

    \I__6617\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34305\
        );

    \I__6616\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34305\
        );

    \I__6615\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34300\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34300\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__34333\,
            I => \N__34297\
        );

    \I__6612\ : CascadeMux
    port map (
            O => \N__34332\,
            I => \N__34293\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__34329\,
            I => \N__34286\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__34326\,
            I => \N__34286\
        );

    \I__6609\ : Span4Mux_h
    port map (
            O => \N__34317\,
            I => \N__34283\
        );

    \I__6608\ : Sp12to4
    port map (
            O => \N__34314\,
            I => \N__34276\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34276\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34300\,
            I => \N__34276\
        );

    \I__6605\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34271\
        );

    \I__6604\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34271\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34264\
        );

    \I__6602\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34264\
        );

    \I__6601\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34264\
        );

    \I__6600\ : Sp12to4
    port map (
            O => \N__34286\,
            I => \N__34261\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__34283\,
            I => \N__34258\
        );

    \I__6598\ : Span12Mux_h
    port map (
            O => \N__34276\,
            I => \N__34251\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__34271\,
            I => \N__34251\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34251\
        );

    \I__6595\ : Odrv12
    port map (
            O => \N__34261\,
            I => n12534
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__34258\,
            I => n12534
        );

    \I__6593\ : Odrv12
    port map (
            O => \N__34251\,
            I => n12534
        );

    \I__6592\ : CascadeMux
    port map (
            O => \N__34244\,
            I => \N__34241\
        );

    \I__6591\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34235\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34235\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34231\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__34234\,
            I => \N__34228\
        );

    \I__6587\ : Span4Mux_v
    port map (
            O => \N__34231\,
            I => \N__34225\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34222\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__34225\,
            I => cmd_rdadctmp_26
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__34222\,
            I => cmd_rdadctmp_26
        );

    \I__6583\ : CEMux
    port map (
            O => \N__34217\,
            I => \N__34213\
        );

    \I__6582\ : CEMux
    port map (
            O => \N__34216\,
            I => \N__34210\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34213\,
            I => \N__34207\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__34210\,
            I => \N__34204\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__34207\,
            I => \N__34201\
        );

    \I__6578\ : Span4Mux_v
    port map (
            O => \N__34204\,
            I => \N__34198\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__34201\,
            I => n12110
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__34198\,
            I => n12110
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__34193\,
            I => \n12110_cascade_\
        );

    \I__6574\ : SRMux
    port map (
            O => \N__34190\,
            I => \N__34186\
        );

    \I__6573\ : SRMux
    port map (
            O => \N__34189\,
            I => \N__34183\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__34186\,
            I => \N__34180\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34177\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__34180\,
            I => \N__34174\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__34177\,
            I => \N__34171\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__34174\,
            I => n14780
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__34171\,
            I => n14780
        );

    \I__6566\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34162\
        );

    \I__6565\ : CascadeMux
    port map (
            O => \N__34165\,
            I => \N__34159\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__34162\,
            I => \N__34156\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34153\
        );

    \I__6562\ : Span4Mux_h
    port map (
            O => \N__34156\,
            I => \N__34150\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__34153\,
            I => data_idxvec_10
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__34150\,
            I => data_idxvec_10
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__34145\,
            I => \n20905_cascade_\
        );

    \I__6558\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34139\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__34139\,
            I => \N__34136\
        );

    \I__6556\ : Span4Mux_v
    port map (
            O => \N__34136\,
            I => \N__34133\
        );

    \I__6555\ : Span4Mux_h
    port map (
            O => \N__34133\,
            I => \N__34130\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__34130\,
            I => n20839
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__34127\,
            I => \n22148_cascade_\
        );

    \I__6552\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34121\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__34121\,
            I => \N__34118\
        );

    \I__6550\ : Span4Mux_h
    port map (
            O => \N__34118\,
            I => \N__34115\
        );

    \I__6549\ : Odrv4
    port map (
            O => \N__34115\,
            I => n22121
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__34112\,
            I => \n22151_cascade_\
        );

    \I__6547\ : CascadeMux
    port map (
            O => \N__34109\,
            I => \n20889_cascade_\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34103\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__34103\,
            I => \N__34100\
        );

    \I__6544\ : Span4Mux_h
    port map (
            O => \N__34100\,
            I => \N__34097\
        );

    \I__6543\ : Span4Mux_h
    port map (
            O => \N__34097\,
            I => \N__34094\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__34094\,
            I => buf_data_iac_18
        );

    \I__6541\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__34088\,
            I => n20906
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \n12152_cascade_\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__6537\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34076\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__34076\,
            I => n12_adj_1639
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__34073\,
            I => \n12194_cascade_\
        );

    \I__6534\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34067\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__34064\,
            I => \N__34060\
        );

    \I__6531\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34057\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__34060\,
            I => \N__34052\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__34057\,
            I => \N__34052\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__34052\,
            I => \N__34048\
        );

    \I__6527\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34045\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__34048\,
            I => \N__34042\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__34045\,
            I => buf_adcdata_iac_0
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__34042\,
            I => buf_adcdata_iac_0
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__34037\,
            I => \n22_cascade_\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34031\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34028\
        );

    \I__6520\ : Span12Mux_h
    port map (
            O => \N__34028\,
            I => \N__34025\
        );

    \I__6519\ : Odrv12
    port map (
            O => \N__34025\,
            I => buf_data_iac_0
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__34022\,
            I => \n30_adj_1484_cascade_\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__34019\,
            I => \N__34016\
        );

    \I__6516\ : InMux
    port map (
            O => \N__34016\,
            I => \N__34013\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__34013\,
            I => \N__34010\
        );

    \I__6514\ : Span4Mux_v
    port map (
            O => \N__34010\,
            I => \N__34007\
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__34007\,
            I => n22_adj_1489
        );

    \I__6512\ : InMux
    port map (
            O => \N__34004\,
            I => \N__34001\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__6510\ : Span4Mux_h
    port map (
            O => \N__33998\,
            I => \N__33995\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__33995\,
            I => \N__33992\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__33992\,
            I => buf_data_iac_1
        );

    \I__6507\ : CascadeMux
    port map (
            O => \N__33989\,
            I => \n30_adj_1504_cascade_\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33983\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__33983\,
            I => \N__33979\
        );

    \I__6504\ : CascadeMux
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__6503\ : Span4Mux_v
    port map (
            O => \N__33979\,
            I => \N__33973\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33970\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__33973\,
            I => buf_adcdata_vdc_0
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33970\,
            I => buf_adcdata_vdc_0
        );

    \I__6499\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33961\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33958\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33954\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33951\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__33957\,
            I => \N__33948\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__33954\,
            I => \N__33945\
        );

    \I__6493\ : Span12Mux_v
    port map (
            O => \N__33951\,
            I => \N__33942\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33939\
        );

    \I__6491\ : Span4Mux_h
    port map (
            O => \N__33945\,
            I => \N__33936\
        );

    \I__6490\ : Span12Mux_h
    port map (
            O => \N__33942\,
            I => \N__33933\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33939\,
            I => buf_adcdata_vac_0
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__33936\,
            I => buf_adcdata_vac_0
        );

    \I__6487\ : Odrv12
    port map (
            O => \N__33933\,
            I => buf_adcdata_vac_0
        );

    \I__6486\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33923\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33923\,
            I => n19_adj_1485
        );

    \I__6484\ : InMux
    port map (
            O => \N__33920\,
            I => \ADC_VDC.genclk.n19494\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33917\,
            I => \ADC_VDC.genclk.n19495\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33914\,
            I => \ADC_VDC.genclk.n19496\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33911\,
            I => \ADC_VDC.genclk.n19497\
        );

    \I__6480\ : CEMux
    port map (
            O => \N__33908\,
            I => \N__33904\
        );

    \I__6479\ : CEMux
    port map (
            O => \N__33907\,
            I => \N__33901\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33898\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33901\,
            I => \N__33895\
        );

    \I__6476\ : Span4Mux_v
    port map (
            O => \N__33898\,
            I => \N__33892\
        );

    \I__6475\ : Span4Mux_v
    port map (
            O => \N__33895\,
            I => \N__33889\
        );

    \I__6474\ : Span4Mux_h
    port map (
            O => \N__33892\,
            I => \N__33886\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__33889\,
            I => \ADC_VDC.genclk.div_state_1__N_1275\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__33886\,
            I => \ADC_VDC.genclk.div_state_1__N_1275\
        );

    \I__6471\ : SRMux
    port map (
            O => \N__33881\,
            I => \N__33877\
        );

    \I__6470\ : SRMux
    port map (
            O => \N__33880\,
            I => \N__33874\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33869\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33866\
        );

    \I__6467\ : SRMux
    port map (
            O => \N__33873\,
            I => \N__33863\
        );

    \I__6466\ : SRMux
    port map (
            O => \N__33872\,
            I => \N__33860\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__33869\,
            I => \N__33857\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__33866\,
            I => \N__33850\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__33863\,
            I => \N__33850\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33850\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__33857\,
            I => \ADC_VDC.genclk.n15067\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__33850\,
            I => \ADC_VDC.genclk.n15067\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33841\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33837\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__33841\,
            I => \N__33834\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33831\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33824\
        );

    \I__6454\ : Span4Mux_v
    port map (
            O => \N__33834\,
            I => \N__33824\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__33831\,
            I => \N__33824\
        );

    \I__6452\ : Span4Mux_h
    port map (
            O => \N__33824\,
            I => \N__33820\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33817\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__33820\,
            I => \N__33814\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__33817\,
            I => \RTD.bit_cnt_3\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__33814\,
            I => \RTD.bit_cnt_3\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33799\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33808\,
            I => \N__33799\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33799\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33796\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33799\,
            I => \RTD.bit_cnt_1\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33796\,
            I => \RTD.bit_cnt_1\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33784\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33784\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33781\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33784\,
            I => \RTD.bit_cnt_2\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33781\,
            I => \RTD.bit_cnt_2\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33772\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__33775\,
            I => \N__33769\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33757\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33757\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33757\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33757\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33754\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__33757\,
            I => \RTD.bit_cnt_0\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__33754\,
            I => \RTD.bit_cnt_0\
        );

    \I__6427\ : CEMux
    port map (
            O => \N__33749\,
            I => \N__33746\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__33743\,
            I => \N__33740\
        );

    \I__6424\ : Span4Mux_h
    port map (
            O => \N__33740\,
            I => \N__33737\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__33737\,
            I => \N__33734\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__33734\,
            I => \RTD.n11756\
        );

    \I__6421\ : SRMux
    port map (
            O => \N__33731\,
            I => \N__33728\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__33725\,
            I => \N__33722\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__6417\ : Span4Mux_h
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6416\ : Odrv4
    port map (
            O => \N__33716\,
            I => \RTD.n15081\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33713\,
            I => \ADC_VDC.genclk.n19485\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33710\,
            I => \ADC_VDC.genclk.n19486\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33707\,
            I => \ADC_VDC.genclk.n19487\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33704\,
            I => \ADC_VDC.genclk.n19488\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33701\,
            I => \ADC_VDC.genclk.n19489\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33698\,
            I => \bfn_13_6_0_\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33695\,
            I => \ADC_VDC.genclk.n19491\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33692\,
            I => \ADC_VDC.genclk.n19492\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33689\,
            I => \ADC_VDC.genclk.n19493\
        );

    \I__6406\ : CEMux
    port map (
            O => \N__33686\,
            I => \N__33683\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33680\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__33680\,
            I => \ADC_VDC.genclk.n6\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33674\,
            I => \N__33670\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33664\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__33670\,
            I => \N__33661\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33654\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33654\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33654\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33664\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__33661\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__33654\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6393\ : CEMux
    port map (
            O => \N__33647\,
            I => \N__33644\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33641\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__33638\,
            I => \N__33635\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__33635\,
            I => \ADC_VDC.n11766\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__33632\,
            I => \N__33625\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__33631\,
            I => \N__33622\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33618\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__33629\,
            I => \N__33615\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33603\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33603\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33603\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33603\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__33618\,
            I => \N__33600\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33597\
        );

    \I__6378\ : CascadeMux
    port map (
            O => \N__33614\,
            I => \N__33594\
        );

    \I__6377\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33589\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33589\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33603\,
            I => \N__33585\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__33600\,
            I => \N__33582\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33579\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33576\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33573\
        );

    \I__6370\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33570\
        );

    \I__6369\ : Span4Mux_v
    port map (
            O => \N__33585\,
            I => \N__33567\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__33582\,
            I => \N__33560\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__33579\,
            I => \N__33560\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__33576\,
            I => \N__33560\
        );

    \I__6365\ : Span4Mux_v
    port map (
            O => \N__33573\,
            I => \N__33555\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33555\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__33567\,
            I => \N__33552\
        );

    \I__6362\ : Span4Mux_v
    port map (
            O => \N__33560\,
            I => \N__33549\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__33555\,
            I => \N__33546\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__33552\,
            I => \N__33543\
        );

    \I__6359\ : Span4Mux_h
    port map (
            O => \N__33549\,
            I => \N__33540\
        );

    \I__6358\ : Span4Mux_h
    port map (
            O => \N__33546\,
            I => \N__33537\
        );

    \I__6357\ : Sp12to4
    port map (
            O => \N__33543\,
            I => \N__33532\
        );

    \I__6356\ : Sp12to4
    port map (
            O => \N__33540\,
            I => \N__33532\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__33537\,
            I => \N__33529\
        );

    \I__6354\ : Odrv12
    port map (
            O => \N__33532\,
            I => \VDC_SDO\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__33529\,
            I => \VDC_SDO\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33511\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33508\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33505\
        );

    \I__6349\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33502\
        );

    \I__6348\ : CascadeMux
    port map (
            O => \N__33520\,
            I => \N__33499\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33494\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33494\
        );

    \I__6345\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33488\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33481\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33481\
        );

    \I__6342\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33481\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__33511\,
            I => \N__33478\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__33508\,
            I => \N__33468\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33465\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33462\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33459\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33494\,
            I => \N__33456\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33451\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33451\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33448\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33488\,
            I => \N__33443\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33481\,
            I => \N__33443\
        );

    \I__6330\ : Span4Mux_h
    port map (
            O => \N__33478\,
            I => \N__33440\
        );

    \I__6329\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33437\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33432\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33432\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33429\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33426\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33421\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33421\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__33468\,
            I => \N__33412\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__33465\,
            I => \N__33412\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__33462\,
            I => \N__33412\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__33459\,
            I => \N__33412\
        );

    \I__6318\ : Span4Mux_h
    port map (
            O => \N__33456\,
            I => \N__33409\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33400\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33448\,
            I => \N__33400\
        );

    \I__6315\ : Span4Mux_h
    port map (
            O => \N__33443\,
            I => \N__33400\
        );

    \I__6314\ : Span4Mux_h
    port map (
            O => \N__33440\,
            I => \N__33400\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__33437\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33432\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33429\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__33426\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__33421\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__33412\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__33409\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__33400\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__33383\,
            I => \N__33380\
        );

    \I__6304\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__33377\,
            I => \ADC_VDC.n62\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__33374\,
            I => \N__33368\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__33373\,
            I => \N__33359\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33355\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__33371\,
            I => \N__33351\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33341\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33322\
        );

    \I__6296\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33322\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33322\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33322\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33322\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33322\
        );

    \I__6291\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33322\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__33358\,
            I => \N__33319\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__33355\,
            I => \N__33316\
        );

    \I__6288\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33311\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33351\,
            I => \N__33311\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33302\
        );

    \I__6285\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33302\
        );

    \I__6284\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33302\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33302\
        );

    \I__6282\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33286\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33286\
        );

    \I__6280\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33280\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33277\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__33340\,
            I => \N__33274\
        );

    \I__6277\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33267\
        );

    \I__6276\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33262\
        );

    \I__6275\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33262\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33259\
        );

    \I__6273\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33256\
        );

    \I__6272\ : Span4Mux_h
    port map (
            O => \N__33316\,
            I => \N__33249\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33249\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33249\
        );

    \I__6269\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33246\
        );

    \I__6268\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33241\
        );

    \I__6267\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33241\
        );

    \I__6266\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33217\
        );

    \I__6265\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33217\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33217\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33217\
        );

    \I__6262\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33217\
        );

    \I__6261\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33217\
        );

    \I__6260\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33217\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33217\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33286\,
            I => \N__33214\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33207\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33207\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33207\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__33280\,
            I => \N__33202\
        );

    \I__6253\ : Span4Mux_v
    port map (
            O => \N__33277\,
            I => \N__33202\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33191\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33191\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33191\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33191\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33191\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__33267\,
            I => \N__33180\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__33262\,
            I => \N__33180\
        );

    \I__6245\ : Span4Mux_h
    port map (
            O => \N__33259\,
            I => \N__33180\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__33256\,
            I => \N__33180\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__33249\,
            I => \N__33180\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33175\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33175\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33172\
        );

    \I__6239\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33167\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33167\
        );

    \I__6237\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33164\
        );

    \I__6236\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33157\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33157\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33157\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33217\,
            I => \N__33146\
        );

    \I__6232\ : Span4Mux_h
    port map (
            O => \N__33214\,
            I => \N__33146\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__33207\,
            I => \N__33146\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__33202\,
            I => \N__33146\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33146\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__33180\,
            I => \N__33141\
        );

    \I__6227\ : Span4Mux_h
    port map (
            O => \N__33175\,
            I => \N__33141\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__33172\,
            I => adc_state_2
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__33167\,
            I => adc_state_2
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__33164\,
            I => adc_state_2
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33157\,
            I => adc_state_2
        );

    \I__6222\ : Odrv4
    port map (
            O => \N__33146\,
            I => adc_state_2
        );

    \I__6221\ : Odrv4
    port map (
            O => \N__33141\,
            I => adc_state_2
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__33128\,
            I => \N__33105\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__33127\,
            I => \N__33102\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__33126\,
            I => \N__33093\
        );

    \I__6217\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33090\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__33124\,
            I => \N__33087\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33076\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33076\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33063\
        );

    \I__6212\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33063\
        );

    \I__6211\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33063\
        );

    \I__6210\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33063\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33063\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33063\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33046\
        );

    \I__6206\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33046\
        );

    \I__6205\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33046\
        );

    \I__6204\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33046\
        );

    \I__6203\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33046\
        );

    \I__6202\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33046\
        );

    \I__6201\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33046\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33046\
        );

    \I__6199\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33035\
        );

    \I__6198\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33035\
        );

    \I__6197\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33035\
        );

    \I__6196\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33028\
        );

    \I__6195\ : InMux
    port map (
            O => \N__33099\,
            I => \N__33028\
        );

    \I__6194\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33028\
        );

    \I__6193\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33023\
        );

    \I__6192\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33023\
        );

    \I__6191\ : InMux
    port map (
            O => \N__33093\,
            I => \N__33019\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__33016\
        );

    \I__6189\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33013\
        );

    \I__6188\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33008\
        );

    \I__6187\ : InMux
    port map (
            O => \N__33085\,
            I => \N__32997\
        );

    \I__6186\ : InMux
    port map (
            O => \N__33084\,
            I => \N__32997\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33083\,
            I => \N__32997\
        );

    \I__6184\ : InMux
    port map (
            O => \N__33082\,
            I => \N__32997\
        );

    \I__6183\ : InMux
    port map (
            O => \N__33081\,
            I => \N__32997\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__32994\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__33063\,
            I => \N__32989\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__32989\
        );

    \I__6179\ : InMux
    port map (
            O => \N__33045\,
            I => \N__32974\
        );

    \I__6178\ : InMux
    port map (
            O => \N__33044\,
            I => \N__32974\
        );

    \I__6177\ : InMux
    port map (
            O => \N__33043\,
            I => \N__32974\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33042\,
            I => \N__32974\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__33035\,
            I => \N__32967\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__32967\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__33023\,
            I => \N__32967\
        );

    \I__6172\ : InMux
    port map (
            O => \N__33022\,
            I => \N__32964\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__32961\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__33016\,
            I => \N__32956\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__33013\,
            I => \N__32956\
        );

    \I__6168\ : InMux
    port map (
            O => \N__33012\,
            I => \N__32951\
        );

    \I__6167\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32951\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__33008\,
            I => \N__32942\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__32997\,
            I => \N__32942\
        );

    \I__6164\ : Span4Mux_v
    port map (
            O => \N__32994\,
            I => \N__32942\
        );

    \I__6163\ : Span4Mux_v
    port map (
            O => \N__32989\,
            I => \N__32942\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32929\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32929\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32929\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32929\
        );

    \I__6158\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32929\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32929\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32924\
        );

    \I__6155\ : Span12Mux_h
    port map (
            O => \N__32967\,
            I => \N__32924\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32964\,
            I => adc_state_3
        );

    \I__6153\ : Odrv4
    port map (
            O => \N__32961\,
            I => adc_state_3
        );

    \I__6152\ : Odrv4
    port map (
            O => \N__32956\,
            I => adc_state_3
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32951\,
            I => adc_state_3
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__32942\,
            I => adc_state_3
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32929\,
            I => adc_state_3
        );

    \I__6148\ : Odrv12
    port map (
            O => \N__32924\,
            I => adc_state_3
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__32909\,
            I => \ADC_VDC.n62_cascade_\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__32906\,
            I => \N__32899\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32887\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32887\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32887\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32884\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32879\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32879\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32876\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32873\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32861\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32861\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32887\,
            I => \N__32852\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__32884\,
            I => \N__32852\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32879\,
            I => \N__32847\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32847\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32842\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32835\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32835\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32835\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32832\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32829\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32824\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32824\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__32861\,
            I => \N__32821\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32818\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32815\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32810\
        );

    \I__6119\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32810\
        );

    \I__6118\ : Span4Mux_h
    port map (
            O => \N__32852\,
            I => \N__32807\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__32847\,
            I => \N__32804\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32799\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32799\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__32842\,
            I => \N__32794\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32794\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32832\,
            I => \N__32785\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32785\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32824\,
            I => \N__32785\
        );

    \I__6109\ : Span12Mux_v
    port map (
            O => \N__32821\,
            I => \N__32785\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32818\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32815\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32810\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6105\ : Odrv4
    port map (
            O => \N__32807\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__32804\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__32799\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__32794\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6101\ : Odrv12
    port map (
            O => \N__32785\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6100\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32765\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32762\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__32762\,
            I => \N__32759\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__32756\,
            I => \ADC_VDC.n11\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32753\,
            I => \bfn_13_5_0_\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32750\,
            I => \ADC_VDC.genclk.n19483\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32747\,
            I => \ADC_VDC.genclk.n19484\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32744\,
            I => n19383
        );

    \I__6091\ : IoInMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__6089\ : Span12Mux_s7_v
    port map (
            O => \N__32735\,
            I => \N__32730\
        );

    \I__6088\ : ClkMux
    port map (
            O => \N__32734\,
            I => \N__32727\
        );

    \I__6087\ : ClkMux
    port map (
            O => \N__32733\,
            I => \N__32724\
        );

    \I__6086\ : Span12Mux_v
    port map (
            O => \N__32730\,
            I => \N__32721\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32718\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32715\
        );

    \I__6083\ : Span12Mux_h
    port map (
            O => \N__32721\,
            I => \N__32711\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__32718\,
            I => \N__32708\
        );

    \I__6081\ : Span4Mux_h
    port map (
            O => \N__32715\,
            I => \N__32705\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32702\
        );

    \I__6079\ : Odrv12
    port map (
            O => \N__32711\,
            I => \TEST_LED\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__32708\,
            I => \TEST_LED\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__32705\,
            I => \TEST_LED\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__32702\,
            I => \TEST_LED\
        );

    \I__6075\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32686\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32683\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32686\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__32683\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__6070\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32674\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32671\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__32674\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32671\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__32666\,
            I => \N__32662\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32659\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__32659\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__32656\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32647\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32644\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32647\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32644\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32636\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__32636\,
            I => \N__32633\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__32633\,
            I => \ADC_VDC.genclk.n27\
        );

    \I__6054\ : CascadeMux
    port map (
            O => \N__32630\,
            I => \ADC_VDC.genclk.n26_cascade_\
        );

    \I__6053\ : CascadeMux
    port map (
            O => \N__32627\,
            I => \ADC_VDC.genclk.n21206_cascade_\
        );

    \I__6052\ : CascadeMux
    port map (
            O => \N__32624\,
            I => \N__32621\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32617\
        );

    \I__6050\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32614\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32617\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__32614\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__6047\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32605\
        );

    \I__6046\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32602\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__32605\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32602\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__6043\ : CascadeMux
    port map (
            O => \N__32597\,
            I => \N__32593\
        );

    \I__6042\ : CascadeMux
    port map (
            O => \N__32596\,
            I => \N__32590\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32587\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32584\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32587\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__32584\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32575\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32572\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__32575\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__32572\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32564\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32564\,
            I => \ADC_VDC.genclk.n21208\
        );

    \I__6031\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32557\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32554\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32557\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__32554\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__32549\,
            I => \N__32546\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32542\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32539\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32542\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__32539\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__32534\,
            I => \N__32530\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32533\,
            I => \N__32527\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32530\,
            I => \N__32524\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__32527\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__32524\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32516\,
            I => \N__32512\
        );

    \I__6015\ : InMux
    port map (
            O => \N__32515\,
            I => \N__32509\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__32512\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__32509\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32501\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__32501\,
            I => \ADC_VDC.genclk.n28\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32495\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__32495\,
            I => \ADC_VDC.genclk.n21206\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32492\,
            I => n19375
        );

    \I__6007\ : InMux
    port map (
            O => \N__32489\,
            I => n19376
        );

    \I__6006\ : InMux
    port map (
            O => \N__32486\,
            I => \bfn_12_18_0_\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32479\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32476\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__32479\,
            I => \N__32473\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__32476\,
            I => acadc_skipcnt_10
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__32473\,
            I => acadc_skipcnt_10
        );

    \I__6000\ : InMux
    port map (
            O => \N__32468\,
            I => n19378
        );

    \I__5999\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32461\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32458\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32455\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__32458\,
            I => acadc_skipcnt_11
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__32455\,
            I => acadc_skipcnt_11
        );

    \I__5994\ : InMux
    port map (
            O => \N__32450\,
            I => n19379
        );

    \I__5993\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32443\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32440\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32437\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__32440\,
            I => acadc_skipcnt_12
        );

    \I__5989\ : Odrv4
    port map (
            O => \N__32437\,
            I => acadc_skipcnt_12
        );

    \I__5988\ : InMux
    port map (
            O => \N__32432\,
            I => n19380
        );

    \I__5987\ : InMux
    port map (
            O => \N__32429\,
            I => n19381
        );

    \I__5986\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32422\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32419\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__32422\,
            I => \N__32416\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32419\,
            I => acadc_skipcnt_14
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__32416\,
            I => acadc_skipcnt_14
        );

    \I__5981\ : InMux
    port map (
            O => \N__32411\,
            I => n19382
        );

    \I__5980\ : InMux
    port map (
            O => \N__32408\,
            I => \bfn_12_17_0_\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32405\,
            I => n19370
        );

    \I__5978\ : InMux
    port map (
            O => \N__32402\,
            I => n19371
        );

    \I__5977\ : InMux
    port map (
            O => \N__32399\,
            I => n19372
        );

    \I__5976\ : InMux
    port map (
            O => \N__32396\,
            I => n19373
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__32393\,
            I => \N__32390\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32386\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32383\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32380\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__32383\,
            I => acadc_skipcnt_6
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__32380\,
            I => acadc_skipcnt_6
        );

    \I__5969\ : InMux
    port map (
            O => \N__32375\,
            I => n19374
        );

    \I__5968\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32368\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__32371\,
            I => \N__32365\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32362\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32358\
        );

    \I__5964\ : Span12Mux_v
    port map (
            O => \N__32362\,
            I => \N__32355\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32352\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__32358\,
            I => \acadc_skipCount_14\
        );

    \I__5961\ : Odrv12
    port map (
            O => \N__32355\,
            I => \acadc_skipCount_14\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__32352\,
            I => \acadc_skipCount_14\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32342\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32334\
        );

    \I__5956\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32329\
        );

    \I__5955\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32329\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__32334\,
            I => \acadc_skipCount_10\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32329\,
            I => \acadc_skipCount_10\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32317\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32314\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__32317\,
            I => acadc_skipcnt_0
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32314\,
            I => acadc_skipcnt_0
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__32309\,
            I => \n16594_cascade_\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32303\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32303\,
            I => n22196
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__32300\,
            I => \n16602_cascade_\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__32294\,
            I => n16602
        );

    \I__5941\ : InMux
    port map (
            O => \N__32291\,
            I => n19407
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__32288\,
            I => \n22169_cascade_\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32282\,
            I => \N__32279\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__5936\ : Span4Mux_v
    port map (
            O => \N__32276\,
            I => \N__32273\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__32273\,
            I => n22079
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__32270\,
            I => \n20568_cascade_\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32263\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32260\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__32263\,
            I => data_idxvec_15
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32260\,
            I => data_idxvec_15
        );

    \I__5929\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32251\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32248\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32251\,
            I => eis_end
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32248\,
            I => eis_end
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__32243\,
            I => \n26_adj_1528_cascade_\
        );

    \I__5924\ : InMux
    port map (
            O => \N__32240\,
            I => \N__32237\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__32237\,
            I => n22166
        );

    \I__5922\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32231\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32231\,
            I => n20742
        );

    \I__5920\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32221\
        );

    \I__5919\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32221\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32218\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__32221\,
            I => \N__32214\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__32217\,
            I => \N__32207\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__32214\,
            I => \N__32204\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32201\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__32210\,
            I => \N__32198\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32195\
        );

    \I__5910\ : Span4Mux_h
    port map (
            O => \N__32204\,
            I => \N__32192\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32189\
        );

    \I__5908\ : Span4Mux_h
    port map (
            O => \N__32198\,
            I => \N__32186\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__32195\,
            I => \N__32181\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__32192\,
            I => \N__32181\
        );

    \I__5905\ : Odrv12
    port map (
            O => \N__32189\,
            I => acadc_trig
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__32186\,
            I => acadc_trig
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__32181\,
            I => acadc_trig
        );

    \I__5902\ : InMux
    port map (
            O => \N__32174\,
            I => n19398
        );

    \I__5901\ : InMux
    port map (
            O => \N__32171\,
            I => n19399
        );

    \I__5900\ : InMux
    port map (
            O => \N__32168\,
            I => \bfn_12_12_0_\
        );

    \I__5899\ : InMux
    port map (
            O => \N__32165\,
            I => n19401
        );

    \I__5898\ : InMux
    port map (
            O => \N__32162\,
            I => n19402
        );

    \I__5897\ : InMux
    port map (
            O => \N__32159\,
            I => n19403
        );

    \I__5896\ : InMux
    port map (
            O => \N__32156\,
            I => n19404
        );

    \I__5895\ : CascadeMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32146\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__32149\,
            I => \N__32143\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__32146\,
            I => \N__32140\
        );

    \I__5891\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32137\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__32140\,
            I => \N__32134\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32137\,
            I => data_idxvec_13
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__32134\,
            I => data_idxvec_13
        );

    \I__5887\ : InMux
    port map (
            O => \N__32129\,
            I => n19405
        );

    \I__5886\ : InMux
    port map (
            O => \N__32126\,
            I => n19406
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__32123\,
            I => \N__32117\
        );

    \I__5884\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32113\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32110\
        );

    \I__5882\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32105\
        );

    \I__5881\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32105\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__32116\,
            I => \N__32102\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32096\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32091\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32091\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32086\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32086\
        );

    \I__5874\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32083\
        );

    \I__5873\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32080\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__32096\,
            I => \N__32077\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__32091\,
            I => \N__32074\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32071\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__32083\,
            I => \N__32068\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__32080\,
            I => \N__32065\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__32077\,
            I => n14522
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__32074\,
            I => n14522
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__32071\,
            I => n14522
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__32068\,
            I => n14522
        );

    \I__5863\ : Odrv12
    port map (
            O => \N__32065\,
            I => n14522
        );

    \I__5862\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32050\
        );

    \I__5861\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32047\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__32041\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32038\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32033\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32033\
        );

    \I__5856\ : CascadeMux
    port map (
            O => \N__32044\,
            I => \N__32029\
        );

    \I__5855\ : Span4Mux_v
    port map (
            O => \N__32041\,
            I => \N__32020\
        );

    \I__5854\ : Span4Mux_h
    port map (
            O => \N__32038\,
            I => \N__32020\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__32033\,
            I => \N__32020\
        );

    \I__5852\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32013\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32029\,
            I => \N__32013\
        );

    \I__5850\ : InMux
    port map (
            O => \N__32028\,
            I => \N__32013\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32010\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__32020\,
            I => n11918
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__32013\,
            I => n11918
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__32010\,
            I => n11918
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__32003\,
            I => \N__31998\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31995\
        );

    \I__5843\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31990\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31990\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__31995\,
            I => cmd_rdadctmp_22
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__31990\,
            I => cmd_rdadctmp_22
        );

    \I__5839\ : InMux
    port map (
            O => \N__31985\,
            I => \bfn_12_11_0_\
        );

    \I__5838\ : InMux
    port map (
            O => \N__31982\,
            I => n19393
        );

    \I__5837\ : InMux
    port map (
            O => \N__31979\,
            I => n19394
        );

    \I__5836\ : InMux
    port map (
            O => \N__31976\,
            I => n19395
        );

    \I__5835\ : InMux
    port map (
            O => \N__31973\,
            I => n19396
        );

    \I__5834\ : InMux
    port map (
            O => \N__31970\,
            I => n19397
        );

    \I__5833\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31962\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31959\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__31965\,
            I => \N__31956\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31962\,
            I => \N__31953\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31959\,
            I => \N__31950\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31947\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__31953\,
            I => \N__31944\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__31950\,
            I => \N__31941\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31947\,
            I => \N__31936\
        );

    \I__5824\ : Sp12to4
    port map (
            O => \N__31944\,
            I => \N__31936\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__31941\,
            I => \N__31933\
        );

    \I__5822\ : Odrv12
    port map (
            O => \N__31936\,
            I => buf_adcdata_vac_22
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__31933\,
            I => buf_adcdata_vac_22
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__31928\,
            I => \N__31925\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31921\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31918\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31921\,
            I => buf_adcdata_vdc_22
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31918\,
            I => buf_adcdata_vdc_22
        );

    \I__5815\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31910\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31910\,
            I => \N__31907\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__31907\,
            I => n22160
        );

    \I__5812\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31900\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31897\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31894\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31897\,
            I => comm_buf_6_4
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__31894\,
            I => comm_buf_6_4
        );

    \I__5807\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31886\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31874\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31869\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31869\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__31877\,
            I => n20646
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__31874\,
            I => n20646
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__31869\,
            I => n20646
        );

    \I__5798\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31859\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31856\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__31856\,
            I => \N__31853\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__31853\,
            I => n30_adj_1630
        );

    \I__5794\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31847\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31844\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__31841\,
            I => n30_adj_1634
        );

    \I__5790\ : InMux
    port map (
            O => \N__31838\,
            I => \N__31835\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31832\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__31829\,
            I => \N__31826\
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__31826\,
            I => n30_adj_1638
        );

    \I__5785\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31820\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31820\,
            I => comm_buf_2_4
        );

    \I__5783\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31814\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__31808\,
            I => n30_adj_1644
        );

    \I__5779\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31802\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__31799\,
            I => \N__31796\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__31796\,
            I => n30_adj_1648
        );

    \I__5775\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31790\,
            I => \N__31786\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__31789\,
            I => \N__31783\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__31786\,
            I => \N__31779\
        );

    \I__5771\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31776\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31773\
        );

    \I__5769\ : Sp12to4
    port map (
            O => \N__31779\,
            I => \N__31768\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__31776\,
            I => \N__31768\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31773\,
            I => cmd_rdadctmp_22_adj_1457
        );

    \I__5766\ : Odrv12
    port map (
            O => \N__31768\,
            I => cmd_rdadctmp_22_adj_1457
        );

    \I__5765\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31760\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__31760\,
            I => \N__31757\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__31757\,
            I => \N__31754\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__31754\,
            I => \ADC_VDC.n10552\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__31751\,
            I => \N__31748\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31745\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__31745\,
            I => \N__31741\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__31744\,
            I => \N__31738\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__31741\,
            I => \N__31735\
        );

    \I__5756\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31732\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__31735\,
            I => \N__31729\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31732\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__31729\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__5752\ : CEMux
    port map (
            O => \N__31724\,
            I => \N__31721\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__31721\,
            I => \ADC_VDC.n12915\
        );

    \I__5750\ : SRMux
    port map (
            O => \N__31718\,
            I => \N__31715\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31712\
        );

    \I__5748\ : Span4Mux_v
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__5747\ : Span4Mux_h
    port map (
            O => \N__31709\,
            I => \N__31706\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__31706\,
            I => \ADC_VDC.n20392\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31703\,
            I => \N__31698\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31695\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31692\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31689\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31695\,
            I => \N__31684\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__31692\,
            I => \N__31684\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__31689\,
            I => \N__31679\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__31684\,
            I => \N__31679\
        );

    \I__5737\ : Span4Mux_h
    port map (
            O => \N__31679\,
            I => \N__31676\
        );

    \I__5736\ : Odrv4
    port map (
            O => \N__31676\,
            I => \RTD.n17720\
        );

    \I__5735\ : SRMux
    port map (
            O => \N__31673\,
            I => \N__31670\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__31670\,
            I => \N__31666\
        );

    \I__5733\ : SRMux
    port map (
            O => \N__31669\,
            I => \N__31663\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__31666\,
            I => \N__31658\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31658\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__31658\,
            I => n14801
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__31655\,
            I => \n2_adj_1587_cascade_\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31649\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31649\,
            I => comm_buf_5_4
        );

    \I__5726\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31643\,
            I => n21324
        );

    \I__5724\ : CascadeMux
    port map (
            O => \N__31640\,
            I => \n4_adj_1588_cascade_\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31637\,
            I => \N__31634\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31634\,
            I => n22136
        );

    \I__5721\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31628\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__31628\,
            I => n1_adj_1586
        );

    \I__5719\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31622\,
            I => n19006
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__31619\,
            I => \n19006_cascade_\
        );

    \I__5716\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31613\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__5714\ : Span12Mux_h
    port map (
            O => \N__31610\,
            I => \N__31607\
        );

    \I__5713\ : Odrv12
    port map (
            O => \N__31607\,
            I => n30_adj_1627
        );

    \I__5712\ : InMux
    port map (
            O => \N__31604\,
            I => \ADC_VDC.genclk.n19482\
        );

    \I__5711\ : CEMux
    port map (
            O => \N__31601\,
            I => \N__31598\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31594\
        );

    \I__5709\ : CEMux
    port map (
            O => \N__31597\,
            I => \N__31591\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__31594\,
            I => \N__31588\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31591\,
            I => \N__31585\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__31588\,
            I => \N__31580\
        );

    \I__5705\ : Span4Mux_v
    port map (
            O => \N__31585\,
            I => \N__31580\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__31580\,
            I => \ADC_VDC.genclk.n11751\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__31577\,
            I => \n12_adj_1615_cascade_\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__31574\,
            I => \n12236_cascade_\
        );

    \I__5701\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31568\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__31565\,
            I => \N__31562\
        );

    \I__5698\ : Sp12to4
    port map (
            O => \N__31562\,
            I => \N__31559\
        );

    \I__5697\ : Odrv12
    port map (
            O => \N__31559\,
            I => buf_data_vac_0
        );

    \I__5696\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__5694\ : Span4Mux_h
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__5693\ : Span4Mux_h
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__5692\ : Span4Mux_h
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__31541\,
            I => buf_data_vac_1
        );

    \I__5690\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31535\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__5687\ : Sp12to4
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__5686\ : Odrv12
    port map (
            O => \N__31526\,
            I => buf_data_vac_2
        );

    \I__5685\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31520\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31520\,
            I => \N__31517\
        );

    \I__5683\ : Span4Mux_h
    port map (
            O => \N__31517\,
            I => \N__31514\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__31514\,
            I => \N__31511\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__31511\,
            I => buf_data_vac_3
        );

    \I__5680\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31505\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31505\,
            I => \N__31502\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__31502\,
            I => \N__31499\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__31496\,
            I => buf_data_vac_4
        );

    \I__5675\ : CEMux
    port map (
            O => \N__31493\,
            I => \N__31490\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__31490\,
            I => \N__31486\
        );

    \I__5673\ : CEMux
    port map (
            O => \N__31489\,
            I => \N__31483\
        );

    \I__5672\ : Span4Mux_v
    port map (
            O => \N__31486\,
            I => \N__31478\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31478\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__31478\,
            I => n12236
        );

    \I__5669\ : InMux
    port map (
            O => \N__31475\,
            I => \ADC_VDC.genclk.n19473\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__31472\,
            I => \N__31468\
        );

    \I__5667\ : InMux
    port map (
            O => \N__31471\,
            I => \N__31465\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31468\,
            I => \N__31462\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__31465\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__31462\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31457\,
            I => \ADC_VDC.genclk.n19474\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31454\,
            I => \bfn_12_4_0_\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31451\,
            I => \ADC_VDC.genclk.n19476\
        );

    \I__5660\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31444\
        );

    \I__5659\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31441\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__31444\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__31441\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31436\,
            I => \ADC_VDC.genclk.n19477\
        );

    \I__5655\ : InMux
    port map (
            O => \N__31433\,
            I => \ADC_VDC.genclk.n19478\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31426\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31423\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31426\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__31423\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31418\,
            I => \ADC_VDC.genclk.n19479\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31415\,
            I => \ADC_VDC.genclk.n19480\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31412\,
            I => \ADC_VDC.genclk.n19481\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__31403\,
            I => \SIG_DDS.tmp_buf_0\
        );

    \I__5644\ : CEMux
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31394\
        );

    \I__5642\ : Span4Mux_v
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__5641\ : Span4Mux_h
    port map (
            O => \N__31391\,
            I => \N__31386\
        );

    \I__5640\ : CEMux
    port map (
            O => \N__31390\,
            I => \N__31383\
        );

    \I__5639\ : CEMux
    port map (
            O => \N__31389\,
            I => \N__31380\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__31386\,
            I => \SIG_DDS.n12738\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31383\,
            I => \SIG_DDS.n12738\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31380\,
            I => \SIG_DDS.n12738\
        );

    \I__5635\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31370\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31366\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31363\
        );

    \I__5632\ : Span4Mux_h
    port map (
            O => \N__31366\,
            I => \N__31360\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31357\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__31360\,
            I => \N__31354\
        );

    \I__5629\ : Span12Mux_h
    port map (
            O => \N__31357\,
            I => \N__31351\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__31354\,
            I => \EIS_SYNCCLK\
        );

    \I__5627\ : Odrv12
    port map (
            O => \N__31351\,
            I => \EIS_SYNCCLK\
        );

    \I__5626\ : IoInMux
    port map (
            O => \N__31346\,
            I => \N__31343\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__31343\,
            I => \N__31340\
        );

    \I__5624\ : Span4Mux_s3_v
    port map (
            O => \N__31340\,
            I => \N__31337\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__31337\,
            I => \OUT_SYNCCLK\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31334\,
            I => \bfn_12_3_0_\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31331\,
            I => \ADC_VDC.genclk.n19468\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__5619\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31321\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31318\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__31321\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__31318\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__5615\ : InMux
    port map (
            O => \N__31313\,
            I => \ADC_VDC.genclk.n19469\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31310\,
            I => \ADC_VDC.genclk.n19470\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31307\,
            I => \ADC_VDC.genclk.n19471\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31304\,
            I => \ADC_VDC.genclk.n19472\
        );

    \I__5611\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31296\
        );

    \I__5610\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31291\
        );

    \I__5609\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31291\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__31296\,
            I => buf_dds0_6
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__31291\,
            I => buf_dds0_6
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__31286\,
            I => \N__31283\
        );

    \I__5605\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31280\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__31280\,
            I => \N__31277\
        );

    \I__5603\ : Span4Mux_h
    port map (
            O => \N__31277\,
            I => \N__31272\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31267\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31267\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__31272\,
            I => buf_dds1_6
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31267\,
            I => buf_dds1_6
        );

    \I__5598\ : CEMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__31259\,
            I => \N__31256\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__31253\,
            I => n11757
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__31250\,
            I => \N__31246\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31241\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31234\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31245\,
            I => \N__31234\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31234\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__31241\,
            I => wdtick_cnt_0
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__31234\,
            I => wdtick_cnt_0
        );

    \I__5587\ : InMux
    port map (
            O => \N__31229\,
            I => \N__31223\
        );

    \I__5586\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31216\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31216\
        );

    \I__5584\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31216\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31223\,
            I => wdtick_cnt_1
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__31216\,
            I => wdtick_cnt_1
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__5580\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31203\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31198\
        );

    \I__5578\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31198\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__31203\,
            I => wdtick_cnt_2
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__31198\,
            I => wdtick_cnt_2
        );

    \I__5575\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31190\,
            I => \N__31185\
        );

    \I__5573\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31182\
        );

    \I__5572\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31179\
        );

    \I__5571\ : Span12Mux_h
    port map (
            O => \N__31185\,
            I => \N__31174\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31174\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__31179\,
            I => buf_dds0_0
        );

    \I__5568\ : Odrv12
    port map (
            O => \N__31174\,
            I => buf_dds0_0
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__31169\,
            I => \n17411_cascade_\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__5565\ : CascadeBuf
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__31160\,
            I => \N__31157\
        );

    \I__5563\ : CascadeBuf
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__31154\,
            I => \N__31151\
        );

    \I__5561\ : CascadeBuf
    port map (
            O => \N__31151\,
            I => \N__31148\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__5559\ : CascadeBuf
    port map (
            O => \N__31145\,
            I => \N__31142\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__5557\ : CascadeBuf
    port map (
            O => \N__31139\,
            I => \N__31136\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__5555\ : CascadeBuf
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__31130\,
            I => \N__31127\
        );

    \I__5553\ : CascadeBuf
    port map (
            O => \N__31127\,
            I => \N__31124\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__31124\,
            I => \N__31121\
        );

    \I__5551\ : CascadeBuf
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__31118\,
            I => \N__31114\
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__31117\,
            I => \N__31111\
        );

    \I__5548\ : CascadeBuf
    port map (
            O => \N__31114\,
            I => \N__31108\
        );

    \I__5547\ : CascadeBuf
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__31108\,
            I => \N__31102\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__31105\,
            I => \N__31099\
        );

    \I__5544\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31096\
        );

    \I__5543\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31093\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__31090\,
            I => \N__31084\
        );

    \I__5539\ : Span12Mux_s9_h
    port map (
            O => \N__31087\,
            I => \N__31081\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__31084\,
            I => \N__31078\
        );

    \I__5537\ : Span12Mux_v
    port map (
            O => \N__31081\,
            I => \N__31075\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__31078\,
            I => \N__31072\
        );

    \I__5535\ : Odrv12
    port map (
            O => \N__31075\,
            I => \data_index_9_N_216_5\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__31072\,
            I => \data_index_9_N_216_5\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31061\
        );

    \I__5532\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31061\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__31061\,
            I => n17409
        );

    \I__5530\ : InMux
    port map (
            O => \N__31058\,
            I => \N__31055\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__31055\,
            I => n17411
        );

    \I__5528\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31047\
        );

    \I__5527\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31044\
        );

    \I__5526\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31041\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__31047\,
            I => data_index_5
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__31044\,
            I => data_index_5
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__31041\,
            I => data_index_5
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__31034\,
            I => \n8828_cascade_\
        );

    \I__5521\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31026\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31023\
        );

    \I__5519\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31020\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__31026\,
            I => data_index_0
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__31023\,
            I => data_index_0
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31020\,
            I => data_index_0
        );

    \I__5515\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__31006\
        );

    \I__5513\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31003\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__31006\,
            I => \N__31000\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31003\,
            I => n8_adj_1532
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__31000\,
            I => n8_adj_1532
        );

    \I__5509\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30990\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30987\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30990\,
            I => \N__30979\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30979\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30974\
        );

    \I__5503\ : Span4Mux_v
    port map (
            O => \N__30979\,
            I => \N__30974\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__30974\,
            I => buf_dds1_13
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30959\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30959\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30959\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30959\,
            I => cmd_rdadctmp_18
        );

    \I__5496\ : IoInMux
    port map (
            O => \N__30956\,
            I => \N__30953\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__5494\ : Span4Mux_s3_h
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__5493\ : Sp12to4
    port map (
            O => \N__30947\,
            I => \N__30943\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30939\
        );

    \I__5491\ : Span12Mux_v
    port map (
            O => \N__30943\,
            I => \N__30936\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30942\,
            I => \N__30933\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30930\
        );

    \I__5488\ : Odrv12
    port map (
            O => \N__30936\,
            I => \AMPV_POW\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30933\,
            I => \AMPV_POW\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__30930\,
            I => \AMPV_POW\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30917\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30917\,
            I => \N__30914\
        );

    \I__5482\ : Odrv12
    port map (
            O => \N__30914\,
            I => n23_adj_1536
        );

    \I__5481\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30904\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30904\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30901\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30904\,
            I => cmd_rdadctmp_21_adj_1429
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30901\,
            I => cmd_rdadctmp_21_adj_1429
        );

    \I__5476\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30892\
        );

    \I__5475\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30889\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30886\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__30889\,
            I => n7_adj_1531
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__30886\,
            I => n7_adj_1531
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__30881\,
            I => \N__30878\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30873\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__30877\,
            I => \N__30870\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__30876\,
            I => \N__30867\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30873\,
            I => \N__30864\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30859\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30859\
        );

    \I__5464\ : Odrv12
    port map (
            O => \N__30864\,
            I => cmd_rdadctmp_22_adj_1428
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30859\,
            I => cmd_rdadctmp_22_adj_1428
        );

    \I__5462\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30851\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__30851\,
            I => \N__30847\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \N__30844\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__30847\,
            I => \N__30841\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30838\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__30841\,
            I => buf_adcdata_vdc_9
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30838\,
            I => buf_adcdata_vdc_9
        );

    \I__5455\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30830\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30830\,
            I => \N__30827\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__30827\,
            I => \N__30824\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__30824\,
            I => \N__30820\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30817\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30814\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30817\,
            I => \N__30808\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__30814\,
            I => \N__30808\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30805\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__30808\,
            I => buf_adcdata_vac_9
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30805\,
            I => buf_adcdata_vac_9
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__5443\ : CascadeBuf
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__5441\ : CascadeBuf
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__5439\ : CascadeBuf
    port map (
            O => \N__30785\,
            I => \N__30782\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \N__30779\
        );

    \I__5437\ : CascadeBuf
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__30776\,
            I => \N__30773\
        );

    \I__5435\ : CascadeBuf
    port map (
            O => \N__30773\,
            I => \N__30770\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__30770\,
            I => \N__30767\
        );

    \I__5433\ : CascadeBuf
    port map (
            O => \N__30767\,
            I => \N__30764\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__30764\,
            I => \N__30761\
        );

    \I__5431\ : CascadeBuf
    port map (
            O => \N__30761\,
            I => \N__30757\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__30760\,
            I => \N__30754\
        );

    \I__5429\ : CascadeMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__5428\ : CascadeBuf
    port map (
            O => \N__30754\,
            I => \N__30748\
        );

    \I__5427\ : CascadeBuf
    port map (
            O => \N__30751\,
            I => \N__30745\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__30748\,
            I => \N__30742\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__30745\,
            I => \N__30739\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30742\,
            I => \N__30736\
        );

    \I__5423\ : CascadeBuf
    port map (
            O => \N__30739\,
            I => \N__30733\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30736\,
            I => \N__30730\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__30733\,
            I => \N__30727\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__30730\,
            I => \N__30724\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__30724\,
            I => \N__30717\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30714\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30711\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__30717\,
            I => \N__30708\
        );

    \I__5414\ : Span12Mux_h
    port map (
            O => \N__30714\,
            I => \N__30705\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30711\,
            I => data_count_8
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__30708\,
            I => data_count_8
        );

    \I__5411\ : Odrv12
    port map (
            O => \N__30705\,
            I => data_count_8
        );

    \I__5410\ : InMux
    port map (
            O => \N__30698\,
            I => \bfn_11_12_0_\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30695\,
            I => n19353
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__5407\ : CascadeBuf
    port map (
            O => \N__30689\,
            I => \N__30686\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__5405\ : CascadeBuf
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__5403\ : CascadeBuf
    port map (
            O => \N__30677\,
            I => \N__30674\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__5401\ : CascadeBuf
    port map (
            O => \N__30671\,
            I => \N__30668\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__30668\,
            I => \N__30665\
        );

    \I__5399\ : CascadeBuf
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__5397\ : CascadeBuf
    port map (
            O => \N__30659\,
            I => \N__30656\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__30656\,
            I => \N__30653\
        );

    \I__5395\ : CascadeBuf
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__30650\,
            I => \N__30647\
        );

    \I__5393\ : CascadeBuf
    port map (
            O => \N__30647\,
            I => \N__30643\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__30646\,
            I => \N__30640\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__30643\,
            I => \N__30637\
        );

    \I__5390\ : CascadeBuf
    port map (
            O => \N__30640\,
            I => \N__30634\
        );

    \I__5389\ : CascadeBuf
    port map (
            O => \N__30637\,
            I => \N__30631\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__30634\,
            I => \N__30628\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__30631\,
            I => \N__30625\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30622\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30619\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__30622\,
            I => \N__30616\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30619\,
            I => \N__30613\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__30616\,
            I => \N__30610\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__30613\,
            I => \N__30607\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__30610\,
            I => \N__30603\
        );

    \I__5379\ : Sp12to4
    port map (
            O => \N__30607\,
            I => \N__30600\
        );

    \I__5378\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30597\
        );

    \I__5377\ : Sp12to4
    port map (
            O => \N__30603\,
            I => \N__30594\
        );

    \I__5376\ : Span12Mux_h
    port map (
            O => \N__30600\,
            I => \N__30591\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30597\,
            I => data_count_9
        );

    \I__5374\ : Odrv12
    port map (
            O => \N__30594\,
            I => data_count_9
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__30591\,
            I => data_count_9
        );

    \I__5372\ : InMux
    port map (
            O => \N__30584\,
            I => \N__30581\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30581\,
            I => \N__30577\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30573\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__30577\,
            I => \N__30570\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__30576\,
            I => \N__30567\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30564\
        );

    \I__5366\ : Span4Mux_h
    port map (
            O => \N__30570\,
            I => \N__30561\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30558\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__30564\,
            I => \N__30555\
        );

    \I__5363\ : Span4Mux_v
    port map (
            O => \N__30561\,
            I => \N__30552\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__30558\,
            I => cmd_rdadctmp_16
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__30555\,
            I => cmd_rdadctmp_16
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__30552\,
            I => cmd_rdadctmp_16
        );

    \I__5359\ : InMux
    port map (
            O => \N__30545\,
            I => \N__30542\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__30542\,
            I => \N__30539\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__30539\,
            I => \N__30536\
        );

    \I__5356\ : Span4Mux_h
    port map (
            O => \N__30536\,
            I => \N__30532\
        );

    \I__5355\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__30532\,
            I => buf_adcdata_vdc_8
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__30529\,
            I => buf_adcdata_vdc_8
        );

    \I__5352\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30518\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__30518\,
            I => \N__30515\
        );

    \I__5349\ : Sp12to4
    port map (
            O => \N__30515\,
            I => \N__30512\
        );

    \I__5348\ : Span12Mux_h
    port map (
            O => \N__30512\,
            I => \N__30507\
        );

    \I__5347\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30502\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30502\
        );

    \I__5345\ : Odrv12
    port map (
            O => \N__30507\,
            I => buf_adcdata_vac_8
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__30502\,
            I => buf_adcdata_vac_8
        );

    \I__5343\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30494\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__30494\,
            I => \N__30491\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__30491\,
            I => \N__30488\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__30488\,
            I => \N__30485\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__30485\,
            I => \N__30481\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30478\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__30481\,
            I => buf_adcdata_vdc_10
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30478\,
            I => buf_adcdata_vdc_10
        );

    \I__5335\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30470\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__30467\,
            I => \N__30464\
        );

    \I__5332\ : Span4Mux_v
    port map (
            O => \N__30464\,
            I => \N__30461\
        );

    \I__5331\ : Sp12to4
    port map (
            O => \N__30461\,
            I => \N__30456\
        );

    \I__5330\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30451\
        );

    \I__5329\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30451\
        );

    \I__5328\ : Odrv12
    port map (
            O => \N__30456\,
            I => buf_adcdata_vac_10
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30451\,
            I => buf_adcdata_vac_10
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__30446\,
            I => \N__30442\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__30445\,
            I => \N__30439\
        );

    \I__5324\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30434\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30434\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__30434\,
            I => \N__30431\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__30431\,
            I => \N__30427\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__30430\,
            I => \N__30424\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__30427\,
            I => \N__30421\
        );

    \I__5318\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30418\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__30421\,
            I => cmd_rdadctmp_17
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__30418\,
            I => cmd_rdadctmp_17
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__30413\,
            I => \n20590_cascade_\
        );

    \I__5314\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30404\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__30404\,
            I => \N__30401\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__30398\,
            I => \N__30393\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30388\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30388\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__30393\,
            I => buf_adcdata_vac_16
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__30388\,
            I => buf_adcdata_vac_16
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5304\ : CascadeBuf
    port map (
            O => \N__30380\,
            I => \N__30377\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__30377\,
            I => \N__30374\
        );

    \I__5302\ : CascadeBuf
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__5300\ : CascadeBuf
    port map (
            O => \N__30368\,
            I => \N__30365\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5298\ : CascadeBuf
    port map (
            O => \N__30362\,
            I => \N__30359\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__30359\,
            I => \N__30356\
        );

    \I__5296\ : CascadeBuf
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__5294\ : CascadeBuf
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5292\ : CascadeBuf
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__30341\,
            I => \N__30338\
        );

    \I__5290\ : CascadeBuf
    port map (
            O => \N__30338\,
            I => \N__30334\
        );

    \I__5289\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \N__30331\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__30334\,
            I => \N__30328\
        );

    \I__5287\ : CascadeBuf
    port map (
            O => \N__30331\,
            I => \N__30325\
        );

    \I__5286\ : CascadeBuf
    port map (
            O => \N__30328\,
            I => \N__30322\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30319\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30310\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30307\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30310\,
            I => \N__30304\
        );

    \I__5279\ : Span4Mux_v
    port map (
            O => \N__30307\,
            I => \N__30300\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__30304\,
            I => \N__30297\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__30303\,
            I => \N__30294\
        );

    \I__5276\ : Sp12to4
    port map (
            O => \N__30300\,
            I => \N__30291\
        );

    \I__5275\ : Sp12to4
    port map (
            O => \N__30297\,
            I => \N__30288\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30285\
        );

    \I__5273\ : Span12Mux_h
    port map (
            O => \N__30291\,
            I => \N__30280\
        );

    \I__5272\ : Span12Mux_h
    port map (
            O => \N__30288\,
            I => \N__30280\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30285\,
            I => data_count_0
        );

    \I__5270\ : Odrv12
    port map (
            O => \N__30280\,
            I => data_count_0
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__5268\ : CascadeBuf
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__5266\ : CascadeBuf
    port map (
            O => \N__30266\,
            I => \N__30263\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__5264\ : CascadeBuf
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__5262\ : CascadeBuf
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__30251\,
            I => \N__30248\
        );

    \I__5260\ : CascadeBuf
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__30245\,
            I => \N__30242\
        );

    \I__5258\ : CascadeBuf
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__30239\,
            I => \N__30236\
        );

    \I__5256\ : CascadeBuf
    port map (
            O => \N__30236\,
            I => \N__30233\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__30233\,
            I => \N__30230\
        );

    \I__5254\ : CascadeBuf
    port map (
            O => \N__30230\,
            I => \N__30226\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__30229\,
            I => \N__30223\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__30226\,
            I => \N__30220\
        );

    \I__5251\ : CascadeBuf
    port map (
            O => \N__30223\,
            I => \N__30217\
        );

    \I__5250\ : CascadeBuf
    port map (
            O => \N__30220\,
            I => \N__30214\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__30217\,
            I => \N__30211\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \N__30208\
        );

    \I__5247\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30205\
        );

    \I__5246\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30202\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__30205\,
            I => \N__30199\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30196\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__30199\,
            I => \N__30193\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__30196\,
            I => \N__30190\
        );

    \I__5241\ : Sp12to4
    port map (
            O => \N__30193\,
            I => \N__30186\
        );

    \I__5240\ : Sp12to4
    port map (
            O => \N__30190\,
            I => \N__30183\
        );

    \I__5239\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30180\
        );

    \I__5238\ : Span12Mux_v
    port map (
            O => \N__30186\,
            I => \N__30175\
        );

    \I__5237\ : Span12Mux_v
    port map (
            O => \N__30183\,
            I => \N__30175\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__30180\,
            I => data_count_1
        );

    \I__5235\ : Odrv12
    port map (
            O => \N__30175\,
            I => data_count_1
        );

    \I__5234\ : InMux
    port map (
            O => \N__30170\,
            I => n19345
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__5232\ : CascadeBuf
    port map (
            O => \N__30164\,
            I => \N__30161\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__5230\ : CascadeBuf
    port map (
            O => \N__30158\,
            I => \N__30155\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__30155\,
            I => \N__30152\
        );

    \I__5228\ : CascadeBuf
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__5227\ : CascadeMux
    port map (
            O => \N__30149\,
            I => \N__30146\
        );

    \I__5226\ : CascadeBuf
    port map (
            O => \N__30146\,
            I => \N__30143\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5224\ : CascadeBuf
    port map (
            O => \N__30140\,
            I => \N__30137\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5222\ : CascadeBuf
    port map (
            O => \N__30134\,
            I => \N__30131\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__5220\ : CascadeBuf
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__5218\ : CascadeBuf
    port map (
            O => \N__30122\,
            I => \N__30119\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__30119\,
            I => \N__30116\
        );

    \I__5216\ : CascadeBuf
    port map (
            O => \N__30116\,
            I => \N__30112\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__30115\,
            I => \N__30109\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__30112\,
            I => \N__30106\
        );

    \I__5213\ : CascadeBuf
    port map (
            O => \N__30109\,
            I => \N__30103\
        );

    \I__5212\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__30103\,
            I => \N__30097\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30094\
        );

    \I__5209\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30091\
        );

    \I__5208\ : Span4Mux_v
    port map (
            O => \N__30094\,
            I => \N__30088\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30085\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__30088\,
            I => \N__30082\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__30085\,
            I => \N__30079\
        );

    \I__5204\ : Sp12to4
    port map (
            O => \N__30082\,
            I => \N__30076\
        );

    \I__5203\ : Sp12to4
    port map (
            O => \N__30079\,
            I => \N__30072\
        );

    \I__5202\ : Span12Mux_h
    port map (
            O => \N__30076\,
            I => \N__30069\
        );

    \I__5201\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30066\
        );

    \I__5200\ : Span12Mux_h
    port map (
            O => \N__30072\,
            I => \N__30061\
        );

    \I__5199\ : Span12Mux_v
    port map (
            O => \N__30069\,
            I => \N__30061\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__30066\,
            I => data_count_2
        );

    \I__5197\ : Odrv12
    port map (
            O => \N__30061\,
            I => data_count_2
        );

    \I__5196\ : InMux
    port map (
            O => \N__30056\,
            I => n19346
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__30053\,
            I => \N__30050\
        );

    \I__5194\ : CascadeBuf
    port map (
            O => \N__30050\,
            I => \N__30047\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__5192\ : CascadeBuf
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__30041\,
            I => \N__30038\
        );

    \I__5190\ : CascadeBuf
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__5188\ : CascadeBuf
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__30029\,
            I => \N__30026\
        );

    \I__5186\ : CascadeBuf
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__30023\,
            I => \N__30020\
        );

    \I__5184\ : CascadeBuf
    port map (
            O => \N__30020\,
            I => \N__30017\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \N__30014\
        );

    \I__5182\ : CascadeBuf
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__30011\,
            I => \N__30008\
        );

    \I__5180\ : CascadeBuf
    port map (
            O => \N__30008\,
            I => \N__30005\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__30005\,
            I => \N__30002\
        );

    \I__5178\ : CascadeBuf
    port map (
            O => \N__30002\,
            I => \N__29998\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__30001\,
            I => \N__29995\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__29998\,
            I => \N__29992\
        );

    \I__5175\ : CascadeBuf
    port map (
            O => \N__29995\,
            I => \N__29989\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29986\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__29989\,
            I => \N__29983\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__29986\,
            I => \N__29980\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29977\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__29980\,
            I => \N__29974\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__5168\ : Sp12to4
    port map (
            O => \N__29974\,
            I => \N__29967\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29964\
        );

    \I__5166\ : Span12Mux_v
    port map (
            O => \N__29970\,
            I => \N__29961\
        );

    \I__5165\ : Span12Mux_h
    port map (
            O => \N__29967\,
            I => \N__29958\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29964\,
            I => data_count_3
        );

    \I__5163\ : Odrv12
    port map (
            O => \N__29961\,
            I => data_count_3
        );

    \I__5162\ : Odrv12
    port map (
            O => \N__29958\,
            I => data_count_3
        );

    \I__5161\ : InMux
    port map (
            O => \N__29951\,
            I => n19347
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__5159\ : CascadeBuf
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5157\ : CascadeBuf
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__29936\,
            I => \N__29933\
        );

    \I__5155\ : CascadeBuf
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__29930\,
            I => \N__29927\
        );

    \I__5153\ : CascadeBuf
    port map (
            O => \N__29927\,
            I => \N__29924\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__29924\,
            I => \N__29921\
        );

    \I__5151\ : CascadeBuf
    port map (
            O => \N__29921\,
            I => \N__29918\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__29918\,
            I => \N__29915\
        );

    \I__5149\ : CascadeBuf
    port map (
            O => \N__29915\,
            I => \N__29912\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__29912\,
            I => \N__29909\
        );

    \I__5147\ : CascadeBuf
    port map (
            O => \N__29909\,
            I => \N__29906\
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__5145\ : CascadeBuf
    port map (
            O => \N__29903\,
            I => \N__29900\
        );

    \I__5144\ : CascadeMux
    port map (
            O => \N__29900\,
            I => \N__29896\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__29899\,
            I => \N__29893\
        );

    \I__5142\ : CascadeBuf
    port map (
            O => \N__29896\,
            I => \N__29890\
        );

    \I__5141\ : CascadeBuf
    port map (
            O => \N__29893\,
            I => \N__29887\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__29890\,
            I => \N__29884\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29881\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29878\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29875\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29878\,
            I => \N__29872\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29875\,
            I => \N__29869\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__29872\,
            I => \N__29866\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__29869\,
            I => \N__29863\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__29866\,
            I => \N__29860\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__29863\,
            I => \N__29856\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__29860\,
            I => \N__29853\
        );

    \I__5129\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29850\
        );

    \I__5128\ : Span4Mux_h
    port map (
            O => \N__29856\,
            I => \N__29847\
        );

    \I__5127\ : Sp12to4
    port map (
            O => \N__29853\,
            I => \N__29844\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__29850\,
            I => data_count_4
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__29847\,
            I => data_count_4
        );

    \I__5124\ : Odrv12
    port map (
            O => \N__29844\,
            I => data_count_4
        );

    \I__5123\ : InMux
    port map (
            O => \N__29837\,
            I => n19348
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5121\ : CascadeBuf
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__5119\ : CascadeBuf
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__29822\,
            I => \N__29819\
        );

    \I__5117\ : CascadeBuf
    port map (
            O => \N__29819\,
            I => \N__29816\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__29816\,
            I => \N__29813\
        );

    \I__5115\ : CascadeBuf
    port map (
            O => \N__29813\,
            I => \N__29810\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__29810\,
            I => \N__29807\
        );

    \I__5113\ : CascadeBuf
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__5111\ : CascadeBuf
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__29798\,
            I => \N__29795\
        );

    \I__5109\ : CascadeBuf
    port map (
            O => \N__29795\,
            I => \N__29792\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__29792\,
            I => \N__29789\
        );

    \I__5107\ : CascadeBuf
    port map (
            O => \N__29789\,
            I => \N__29786\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__29786\,
            I => \N__29782\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__29785\,
            I => \N__29779\
        );

    \I__5104\ : CascadeBuf
    port map (
            O => \N__29782\,
            I => \N__29776\
        );

    \I__5103\ : CascadeBuf
    port map (
            O => \N__29779\,
            I => \N__29773\
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__29776\,
            I => \N__29770\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__29773\,
            I => \N__29767\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29764\
        );

    \I__5099\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29764\,
            I => \N__29758\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29754\
        );

    \I__5096\ : Sp12to4
    port map (
            O => \N__29758\,
            I => \N__29751\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29748\
        );

    \I__5094\ : Span12Mux_h
    port map (
            O => \N__29754\,
            I => \N__29745\
        );

    \I__5093\ : Span12Mux_v
    port map (
            O => \N__29751\,
            I => \N__29742\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29748\,
            I => data_count_5
        );

    \I__5091\ : Odrv12
    port map (
            O => \N__29745\,
            I => data_count_5
        );

    \I__5090\ : Odrv12
    port map (
            O => \N__29742\,
            I => data_count_5
        );

    \I__5089\ : InMux
    port map (
            O => \N__29735\,
            I => n19349
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__5087\ : CascadeBuf
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__29726\,
            I => \N__29723\
        );

    \I__5085\ : CascadeBuf
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__5083\ : CascadeBuf
    port map (
            O => \N__29717\,
            I => \N__29714\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__5081\ : CascadeBuf
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__29708\,
            I => \N__29705\
        );

    \I__5079\ : CascadeBuf
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__29702\,
            I => \N__29699\
        );

    \I__5077\ : CascadeBuf
    port map (
            O => \N__29699\,
            I => \N__29696\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__29696\,
            I => \N__29693\
        );

    \I__5075\ : CascadeBuf
    port map (
            O => \N__29693\,
            I => \N__29690\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__29690\,
            I => \N__29686\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__29689\,
            I => \N__29683\
        );

    \I__5072\ : CascadeBuf
    port map (
            O => \N__29686\,
            I => \N__29680\
        );

    \I__5071\ : CascadeBuf
    port map (
            O => \N__29683\,
            I => \N__29677\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29674\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__29677\,
            I => \N__29671\
        );

    \I__5068\ : CascadeBuf
    port map (
            O => \N__29674\,
            I => \N__29668\
        );

    \I__5067\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29665\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__29668\,
            I => \N__29662\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29659\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29656\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__29659\,
            I => \N__29653\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29656\,
            I => \N__29650\
        );

    \I__5061\ : Span4Mux_v
    port map (
            O => \N__29653\,
            I => \N__29646\
        );

    \I__5060\ : Sp12to4
    port map (
            O => \N__29650\,
            I => \N__29643\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29640\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__29646\,
            I => \N__29637\
        );

    \I__5057\ : Span12Mux_v
    port map (
            O => \N__29643\,
            I => \N__29634\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29640\,
            I => data_count_6
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__29637\,
            I => data_count_6
        );

    \I__5054\ : Odrv12
    port map (
            O => \N__29634\,
            I => data_count_6
        );

    \I__5053\ : InMux
    port map (
            O => \N__29627\,
            I => n19350
        );

    \I__5052\ : CascadeMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__5051\ : CascadeBuf
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__29618\,
            I => \N__29615\
        );

    \I__5049\ : CascadeBuf
    port map (
            O => \N__29615\,
            I => \N__29612\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__5047\ : CascadeBuf
    port map (
            O => \N__29609\,
            I => \N__29606\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__29606\,
            I => \N__29603\
        );

    \I__5045\ : CascadeBuf
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__29600\,
            I => \N__29597\
        );

    \I__5043\ : CascadeBuf
    port map (
            O => \N__29597\,
            I => \N__29594\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__29594\,
            I => \N__29591\
        );

    \I__5041\ : CascadeBuf
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5039\ : CascadeBuf
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__5037\ : CascadeBuf
    port map (
            O => \N__29579\,
            I => \N__29575\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__29578\,
            I => \N__29572\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__5034\ : CascadeBuf
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__5033\ : CascadeBuf
    port map (
            O => \N__29569\,
            I => \N__29563\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__29563\,
            I => \N__29557\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29554\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29551\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__29554\,
            I => \N__29548\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__29551\,
            I => \N__29545\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__29548\,
            I => \N__29542\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__29545\,
            I => \N__29539\
        );

    \I__5024\ : Sp12to4
    port map (
            O => \N__29542\,
            I => \N__29535\
        );

    \I__5023\ : Sp12to4
    port map (
            O => \N__29539\,
            I => \N__29532\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29529\
        );

    \I__5021\ : Span12Mux_v
    port map (
            O => \N__29535\,
            I => \N__29524\
        );

    \I__5020\ : Span12Mux_v
    port map (
            O => \N__29532\,
            I => \N__29524\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29529\,
            I => data_count_7
        );

    \I__5018\ : Odrv12
    port map (
            O => \N__29524\,
            I => data_count_7
        );

    \I__5017\ : InMux
    port map (
            O => \N__29519\,
            I => n19351
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__29516\,
            I => \N__29512\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__29515\,
            I => \N__29509\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29505\
        );

    \I__5013\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29502\
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__29508\,
            I => \N__29499\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29496\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29492\
        );

    \I__5009\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29489\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__29496\,
            I => \N__29485\
        );

    \I__5007\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29482\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__29492\,
            I => \N__29479\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__29489\,
            I => \N__29476\
        );

    \I__5004\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29473\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__29485\,
            I => \N__29468\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__29482\,
            I => \N__29468\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__29479\,
            I => \buf_cfgRTD_6\
        );

    \I__5000\ : Odrv12
    port map (
            O => \N__29476\,
            I => \buf_cfgRTD_6\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__29473\,
            I => \buf_cfgRTD_6\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__29468\,
            I => \buf_cfgRTD_6\
        );

    \I__4997\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29456\,
            I => \N__29453\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__29453\,
            I => \N__29448\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__29452\,
            I => \N__29445\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__29448\,
            I => \N__29439\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29434\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29434\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__29439\,
            I => cmd_rdadctmp_27
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__29434\,
            I => cmd_rdadctmp_27
        );

    \I__4987\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29425\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29422\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29425\,
            I => \N__29418\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__29422\,
            I => \N__29415\
        );

    \I__4983\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29412\
        );

    \I__4982\ : Span12Mux_h
    port map (
            O => \N__29418\,
            I => \N__29409\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__29415\,
            I => \N__29406\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__29412\,
            I => buf_adcdata_vac_19
        );

    \I__4979\ : Odrv12
    port map (
            O => \N__29409\,
            I => buf_adcdata_vac_19
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__29406\,
            I => buf_adcdata_vac_19
        );

    \I__4977\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29395\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__29398\,
            I => \N__29391\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__29395\,
            I => \N__29388\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \N__29385\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29382\
        );

    \I__4972\ : Span12Mux_h
    port map (
            O => \N__29388\,
            I => \N__29379\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29376\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__29382\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4969\ : Odrv12
    port map (
            O => \N__29379\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__29376\,
            I => cmd_rdadctmp_8_adj_1442
        );

    \I__4967\ : CascadeMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__4966\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29359\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29359\
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__29364\,
            I => \N__29356\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29359\,
            I => \N__29353\
        );

    \I__4962\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29350\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__29353\,
            I => cmd_rdadctmp_9_adj_1441
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__29350\,
            I => cmd_rdadctmp_9_adj_1441
        );

    \I__4959\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29342\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29338\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__29341\,
            I => \N__29335\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__29338\,
            I => \N__29332\
        );

    \I__4955\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29329\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__29332\,
            I => buf_adcdata_vdc_15
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__29329\,
            I => buf_adcdata_vdc_15
        );

    \I__4952\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29318\
        );

    \I__4950\ : Span4Mux_v
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__29315\,
            I => \N__29312\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__29312\,
            I => \N__29307\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29302\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29302\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__29307\,
            I => buf_adcdata_vac_15
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29302\,
            I => buf_adcdata_vac_15
        );

    \I__4943\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29294\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__29288\,
            I => n22016
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__29285\,
            I => \N__29282\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29275\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__29275\,
            I => \N__29269\
        );

    \I__4934\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29266\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__29269\,
            I => buf_adcdata_vdc_16
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29266\,
            I => buf_adcdata_vdc_16
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__29261\,
            I => \N__29257\
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \N__29253\
        );

    \I__4929\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29250\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29245\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29245\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29250\,
            I => cmd_rdadctmp_23
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__29245\,
            I => cmd_rdadctmp_23
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__29240\,
            I => \N__29235\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29232\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29229\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29226\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29223\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__29229\,
            I => cmd_rdadctmp_24
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29226\,
            I => cmd_rdadctmp_24
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__29223\,
            I => cmd_rdadctmp_24
        );

    \I__4916\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29212\
        );

    \I__4915\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29209\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29212\,
            I => cmd_rdadcbuf_27
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29209\,
            I => cmd_rdadcbuf_27
        );

    \I__4912\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29201\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__29201\,
            I => \N__29197\
        );

    \I__4910\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29194\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__29197\,
            I => cmd_rdadcbuf_11
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__29194\,
            I => cmd_rdadcbuf_11
        );

    \I__4907\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29185\
        );

    \I__4906\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29182\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__29185\,
            I => cmd_rdadcbuf_33
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29182\,
            I => cmd_rdadcbuf_33
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29154\
        );

    \I__4901\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29154\
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__29172\,
            I => \N__29151\
        );

    \I__4899\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29147\
        );

    \I__4898\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29132\
        );

    \I__4897\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29132\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29132\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29132\
        );

    \I__4894\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29132\
        );

    \I__4893\ : InMux
    port map (
            O => \N__29165\,
            I => \N__29132\
        );

    \I__4892\ : InMux
    port map (
            O => \N__29164\,
            I => \N__29132\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__29163\,
            I => \N__29128\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__29162\,
            I => \N__29121\
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__29161\,
            I => \N__29118\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__29160\,
            I => \N__29115\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__29159\,
            I => \N__29112\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__29154\,
            I => \N__29107\
        );

    \I__4885\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29102\
        );

    \I__4884\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29102\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29147\,
            I => \N__29099\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__29132\,
            I => \N__29096\
        );

    \I__4881\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29093\
        );

    \I__4880\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29090\
        );

    \I__4879\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29073\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29073\
        );

    \I__4877\ : InMux
    port map (
            O => \N__29125\,
            I => \N__29073\
        );

    \I__4876\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29073\
        );

    \I__4875\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29073\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29073\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29073\
        );

    \I__4872\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29073\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29068\
        );

    \I__4870\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29068\
        );

    \I__4869\ : Span4Mux_v
    port map (
            O => \N__29107\,
            I => \N__29065\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__29102\,
            I => \N__29058\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__29099\,
            I => \N__29058\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__29096\,
            I => \N__29058\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__29093\,
            I => n13109
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__29090\,
            I => n13109
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__29073\,
            I => n13109
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__29068\,
            I => n13109
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__29065\,
            I => n13109
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__29058\,
            I => n13109
        );

    \I__4859\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29041\
        );

    \I__4858\ : InMux
    port map (
            O => \N__29044\,
            I => \N__29038\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__29041\,
            I => cmd_rdadcbuf_20
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__29038\,
            I => cmd_rdadcbuf_20
        );

    \I__4855\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__29030\,
            I => \N__29025\
        );

    \I__4853\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29022\
        );

    \I__4852\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29019\
        );

    \I__4851\ : Span12Mux_h
    port map (
            O => \N__29025\,
            I => \N__29016\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__29013\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__29019\,
            I => buf_adcdata_vac_18
        );

    \I__4848\ : Odrv12
    port map (
            O => \N__29016\,
            I => buf_adcdata_vac_18
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__29013\,
            I => buf_adcdata_vac_18
        );

    \I__4846\ : InMux
    port map (
            O => \N__29006\,
            I => \N__29002\
        );

    \I__4845\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28997\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28991\
        );

    \I__4843\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28986\
        );

    \I__4842\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28986\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28997\,
            I => \N__28983\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28980\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28974\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28974\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28969\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__28986\,
            I => \N__28969\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__28983\,
            I => \N__28964\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28980\,
            I => \N__28964\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28961\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28958\
        );

    \I__4831\ : Span4Mux_v
    port map (
            O => \N__28969\,
            I => \N__28955\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__28964\,
            I => \N__28952\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28947\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__28958\,
            I => \N__28947\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28955\,
            I => n12411
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__28952\,
            I => n12411
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__28947\,
            I => n12411
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__28940\,
            I => \n30_adj_1480_cascade_\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__4820\ : Span4Mux_v
    port map (
            O => \N__28930\,
            I => \N__28924\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__28924\,
            I => buf_adcdata_vdc_1
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28921\,
            I => buf_adcdata_vdc_1
        );

    \I__4816\ : CascadeMux
    port map (
            O => \N__28916\,
            I => \n19_adj_1491_cascade_\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__4813\ : Span12Mux_h
    port map (
            O => \N__28907\,
            I => \N__28902\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28897\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28897\
        );

    \I__4810\ : Odrv12
    port map (
            O => \N__28902\,
            I => buf_adcdata_iac_1
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28897\,
            I => buf_adcdata_iac_1
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__28892\,
            I => \N__28889\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28886\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28882\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28879\
        );

    \I__4804\ : Span4Mux_v
    port map (
            O => \N__28882\,
            I => \N__28874\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28879\,
            I => \N__28874\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__28874\,
            I => \buf_readRTD_14\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28867\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28867\,
            I => cmd_rdadcbuf_26
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__28864\,
            I => cmd_rdadcbuf_26
        );

    \I__4797\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28855\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28852\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28855\,
            I => cmd_rdadcbuf_25
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__28852\,
            I => cmd_rdadcbuf_25
        );

    \I__4793\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28843\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28840\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__28843\,
            I => cmd_rdadcbuf_24
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28840\,
            I => cmd_rdadcbuf_24
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__28835\,
            I => \N__28831\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__28834\,
            I => \N__28828\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28825\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28821\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28818\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__28824\,
            I => \N__28815\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28821\,
            I => \N__28810\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__28818\,
            I => \N__28810\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28807\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__28810\,
            I => cmd_rdadctmp_11
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28807\,
            I => cmd_rdadctmp_11
        );

    \I__4778\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__4776\ : Span12Mux_h
    port map (
            O => \N__28796\,
            I => \N__28791\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28786\
        );

    \I__4774\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28786\
        );

    \I__4773\ : Odrv12
    port map (
            O => \N__28791\,
            I => buf_adcdata_vac_3
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__28786\,
            I => buf_adcdata_vac_3
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__28781\,
            I => \N__28777\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__28780\,
            I => \N__28773\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28766\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28766\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28766\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28766\,
            I => cmd_rdadctmp_11_adj_1439
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__28763\,
            I => \N__28759\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__28762\,
            I => \N__28756\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28752\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28749\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__28755\,
            I => \N__28746\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28743\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__28749\,
            I => \N__28740\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28737\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__28743\,
            I => \N__28734\
        );

    \I__4756\ : Span4Mux_v
    port map (
            O => \N__28740\,
            I => \N__28731\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28737\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__28734\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__28731\,
            I => cmd_rdadctmp_12_adj_1438
        );

    \I__4752\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28721\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__28718\,
            I => \N__28715\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__28715\,
            I => \N__28712\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__28712\,
            I => \N__28709\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__28709\,
            I => buf_data_vac_7
        );

    \I__4746\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28703\,
            I => \N__28700\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__28700\,
            I => \N__28697\
        );

    \I__4743\ : Span4Mux_h
    port map (
            O => \N__28697\,
            I => \N__28694\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__28694\,
            I => buf_data_vac_6
        );

    \I__4741\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28688\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28688\,
            I => \N__28685\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__28685\,
            I => \N__28682\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__28682\,
            I => \N__28679\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__28679\,
            I => buf_data_vac_5
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28670\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28670\,
            I => \N__28665\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28662\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__28668\,
            I => \N__28659\
        );

    \I__4731\ : Span4Mux_v
    port map (
            O => \N__28665\,
            I => \N__28656\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28662\,
            I => \N__28653\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28650\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__28656\,
            I => cmd_rdadctmp_10_adj_1440
        );

    \I__4727\ : Odrv12
    port map (
            O => \N__28653\,
            I => cmd_rdadctmp_10_adj_1440
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28650\,
            I => cmd_rdadctmp_10_adj_1440
        );

    \I__4725\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28640\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28640\,
            I => \N__28637\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__28637\,
            I => \N__28633\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__28636\,
            I => \N__28630\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__28633\,
            I => \N__28627\
        );

    \I__4720\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28624\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28627\,
            I => buf_adcdata_vdc_2
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__28624\,
            I => buf_adcdata_vdc_2
        );

    \I__4717\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__28610\,
            I => \N__28607\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__28607\,
            I => \N__28602\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28597\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28597\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__28602\,
            I => buf_adcdata_vac_2
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__28597\,
            I => buf_adcdata_vac_2
        );

    \I__4708\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28589\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__28586\,
            I => \N__28582\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28578\
        );

    \I__4704\ : Sp12to4
    port map (
            O => \N__28582\,
            I => \N__28575\
        );

    \I__4703\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28572\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28578\,
            I => buf_adcdata_iac_2
        );

    \I__4701\ : Odrv12
    port map (
            O => \N__28575\,
            I => buf_adcdata_iac_2
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__28572\,
            I => buf_adcdata_iac_2
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__28565\,
            I => \n19_adj_1646_cascade_\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28556\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__28556\,
            I => \N__28553\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__28553\,
            I => \N__28550\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__28550\,
            I => \N__28547\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__28547\,
            I => buf_data_iac_2
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__28544\,
            I => \n22_adj_1647_cascade_\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__28541\,
            I => \N__28538\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28532\
        );

    \I__4689\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28532\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28528\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__28531\,
            I => \N__28525\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__28528\,
            I => \N__28522\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28519\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__28522\,
            I => cmd_rdadctmp_10
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__28519\,
            I => cmd_rdadctmp_10
        );

    \I__4682\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28507\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28504\
        );

    \I__4679\ : Span4Mux_v
    port map (
            O => \N__28507\,
            I => \N__28501\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28504\,
            I => \N__28498\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__28501\,
            I => buf_adcdata_vdc_3
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__28498\,
            I => buf_adcdata_vdc_3
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__28493\,
            I => \n19_adj_1642_cascade_\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28487\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__28481\,
            I => \N__28478\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__28478\,
            I => buf_data_iac_3
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__28475\,
            I => \n22_adj_1643_cascade_\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__4666\ : Span12Mux_h
    port map (
            O => \N__28466\,
            I => \N__28461\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28456\
        );

    \I__4664\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28456\
        );

    \I__4663\ : Odrv12
    port map (
            O => \N__28461\,
            I => buf_adcdata_iac_3
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__28456\,
            I => buf_adcdata_iac_3
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__28451\,
            I => \N__28448\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__28445\,
            I => \SIG_DDS.tmp_buf_5\
        );

    \I__4658\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28437\
        );

    \I__4657\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28434\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28431\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28428\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28434\,
            I => buf_dds0_2
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__28431\,
            I => buf_dds0_2
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__28428\,
            I => buf_dds0_2
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__28421\,
            I => \N__28418\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28415\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__28415\,
            I => \N__28410\
        );

    \I__4648\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28407\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28413\,
            I => \N__28404\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__28410\,
            I => \N__28401\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28407\,
            I => \N__28398\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28404\,
            I => buf_dds0_4
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__28401\,
            I => buf_dds0_4
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__28398\,
            I => buf_dds0_4
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__4640\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28385\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28385\,
            I => \SIG_DDS.tmp_buf_4\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4637\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28376\,
            I => \SIG_DDS.tmp_buf_7\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28369\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__28372\,
            I => \N__28365\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__28369\,
            I => \N__28362\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28357\
        );

    \I__4631\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28357\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__28362\,
            I => buf_dds0_8
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28357\,
            I => buf_dds0_8
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__4627\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28346\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28346\,
            I => \N__28343\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__28343\,
            I => \SIG_DDS.tmp_buf_8\
        );

    \I__4624\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28336\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28332\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28329\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28326\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__28332\,
            I => \N__28323\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__28329\,
            I => buf_dds0_1
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28326\,
            I => buf_dds0_1
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__28323\,
            I => buf_dds0_1
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28310\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__28310\,
            I => \SIG_DDS.tmp_buf_1\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__28307\,
            I => \N__28304\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28301\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__28301\,
            I => \SIG_DDS.tmp_buf_2\
        );

    \I__4610\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__4608\ : Span4Mux_h
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__4607\ : Span4Mux_v
    port map (
            O => \N__28289\,
            I => \N__28284\
        );

    \I__4606\ : InMux
    port map (
            O => \N__28288\,
            I => \N__28281\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28278\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__28284\,
            I => buf_dds0_3
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__28281\,
            I => buf_dds0_3
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28278\,
            I => buf_dds0_3
        );

    \I__4601\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__28268\,
            I => \SIG_DDS.tmp_buf_3\
        );

    \I__4599\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__4597\ : Odrv12
    port map (
            O => \N__28259\,
            I => n8_adj_1553
        );

    \I__4596\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28252\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__28249\,
            I => n7_adj_1552
        );

    \I__4592\ : Odrv12
    port map (
            O => \N__28246\,
            I => n7_adj_1552
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__4590\ : CascadeBuf
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__28235\,
            I => \N__28232\
        );

    \I__4588\ : CascadeBuf
    port map (
            O => \N__28232\,
            I => \N__28229\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__4586\ : CascadeBuf
    port map (
            O => \N__28226\,
            I => \N__28223\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__4584\ : CascadeBuf
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__28217\,
            I => \N__28214\
        );

    \I__4582\ : CascadeBuf
    port map (
            O => \N__28214\,
            I => \N__28211\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__28211\,
            I => \N__28208\
        );

    \I__4580\ : CascadeBuf
    port map (
            O => \N__28208\,
            I => \N__28205\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__28205\,
            I => \N__28201\
        );

    \I__4578\ : CascadeMux
    port map (
            O => \N__28204\,
            I => \N__28198\
        );

    \I__4577\ : CascadeBuf
    port map (
            O => \N__28201\,
            I => \N__28195\
        );

    \I__4576\ : CascadeBuf
    port map (
            O => \N__28198\,
            I => \N__28192\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__28195\,
            I => \N__28189\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__28192\,
            I => \N__28186\
        );

    \I__4573\ : CascadeBuf
    port map (
            O => \N__28189\,
            I => \N__28183\
        );

    \I__4572\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28180\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__28183\,
            I => \N__28177\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28174\
        );

    \I__4569\ : CascadeBuf
    port map (
            O => \N__28177\,
            I => \N__28171\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__28174\,
            I => \N__28168\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__28171\,
            I => \N__28165\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__28168\,
            I => \N__28162\
        );

    \I__4565\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28159\
        );

    \I__4564\ : Sp12to4
    port map (
            O => \N__28162\,
            I => \N__28156\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28159\,
            I => \N__28153\
        );

    \I__4562\ : Span12Mux_v
    port map (
            O => \N__28156\,
            I => \N__28148\
        );

    \I__4561\ : Span12Mux_s8_h
    port map (
            O => \N__28153\,
            I => \N__28148\
        );

    \I__4560\ : Odrv12
    port map (
            O => \N__28148\,
            I => \data_index_9_N_216_9\
        );

    \I__4559\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28140\
        );

    \I__4558\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28135\
        );

    \I__4557\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28135\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__28140\,
            I => buf_dds0_10
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28135\,
            I => buf_dds0_10
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__28130\,
            I => \N__28127\
        );

    \I__4553\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28124\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__28124\,
            I => \SIG_DDS.tmp_buf_10\
        );

    \I__4551\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28118\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28113\
        );

    \I__4549\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28110\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28107\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__28113\,
            I => \N__28102\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__28110\,
            I => \N__28102\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__28107\,
            I => buf_dds0_13
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__28102\,
            I => buf_dds0_13
        );

    \I__4543\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__28094\,
            I => \SIG_DDS.tmp_buf_13\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__28088\,
            I => \SIG_DDS.tmp_buf_11\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__28085\,
            I => \N__28082\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4536\ : Odrv12
    port map (
            O => \N__28076\,
            I => \SIG_DDS.tmp_buf_12\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__4534\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__28067\,
            I => \SIG_DDS.tmp_buf_14\
        );

    \I__4532\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28057\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28053\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__28057\,
            I => \N__28050\
        );

    \I__4528\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28047\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28044\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__28050\,
            I => \N__28041\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__28047\,
            I => buf_dds0_15
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__28044\,
            I => buf_dds0_15
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__28041\,
            I => buf_dds0_15
        );

    \I__4522\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__28027\
        );

    \I__4520\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28024\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__28027\,
            I => \N__28020\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__28017\
        );

    \I__4517\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28014\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__28020\,
            I => buf_dds0_9
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__28017\,
            I => buf_dds0_9
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__28014\,
            I => buf_dds0_9
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__4512\ : InMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__28001\,
            I => \SIG_DDS.tmp_buf_9\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27992\,
            I => \SIG_DDS.tmp_buf_6\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__27989\,
            I => \n8_adj_1553_cascade_\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27981\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27976\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27976\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__27981\,
            I => data_index_9
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27976\,
            I => data_index_9
        );

    \I__4501\ : IoInMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__4499\ : IoSpan4Mux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__4498\ : Span4Mux_s2_h
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__4497\ : Span4Mux_h
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__4496\ : Sp12to4
    port map (
            O => \N__27956\,
            I => \N__27953\
        );

    \I__4495\ : Span12Mux_v
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__4494\ : Span12Mux_h
    port map (
            O => \N__27950\,
            I => \N__27947\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__27947\,
            I => \ICE_GPMI_0\
        );

    \I__4492\ : CEMux
    port map (
            O => \N__27944\,
            I => \N__27941\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27938\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__27938\,
            I => n11401
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__27935\,
            I => \n20772_cascade_\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__27932\,
            I => \n11835_cascade_\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27929\,
            I => n19388
        );

    \I__4486\ : InMux
    port map (
            O => \N__27926\,
            I => n19389
        );

    \I__4485\ : InMux
    port map (
            O => \N__27923\,
            I => n19390
        );

    \I__4484\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27916\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27913\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27907\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27913\,
            I => \N__27907\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27904\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__27907\,
            I => data_index_8
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27904\,
            I => data_index_8
        );

    \I__4477\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27893\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27893\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27893\,
            I => n7_adj_1554
        );

    \I__4474\ : InMux
    port map (
            O => \N__27890\,
            I => \bfn_10_15_0_\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27887\,
            I => n19392
        );

    \I__4472\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27880\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27876\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__27880\,
            I => \N__27873\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27870\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27876\,
            I => buf_dds1_2
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__27873\,
            I => buf_dds1_2
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27870\,
            I => buf_dds1_2
        );

    \I__4465\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27858\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27855\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27852\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27858\,
            I => data_index_7
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__27855\,
            I => data_index_7
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__27852\,
            I => data_index_7
        );

    \I__4459\ : InMux
    port map (
            O => \N__27845\,
            I => \N__27842\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27842\,
            I => n8_adj_1557
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \n8_adj_1557_cascade_\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27832\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27829\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27832\,
            I => n7_adj_1556
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27829\,
            I => n7_adj_1556
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__27824\,
            I => \N__27821\
        );

    \I__4451\ : CascadeBuf
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__4449\ : CascadeBuf
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__27812\,
            I => \N__27809\
        );

    \I__4447\ : CascadeBuf
    port map (
            O => \N__27809\,
            I => \N__27806\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__4445\ : CascadeBuf
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__27800\,
            I => \N__27797\
        );

    \I__4443\ : CascadeBuf
    port map (
            O => \N__27797\,
            I => \N__27794\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__27794\,
            I => \N__27791\
        );

    \I__4441\ : CascadeBuf
    port map (
            O => \N__27791\,
            I => \N__27788\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__27788\,
            I => \N__27785\
        );

    \I__4439\ : CascadeBuf
    port map (
            O => \N__27785\,
            I => \N__27782\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__27782\,
            I => \N__27778\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__4436\ : CascadeBuf
    port map (
            O => \N__27778\,
            I => \N__27772\
        );

    \I__4435\ : CascadeBuf
    port map (
            O => \N__27775\,
            I => \N__27769\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__27772\,
            I => \N__27766\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__27769\,
            I => \N__27763\
        );

    \I__4432\ : CascadeBuf
    port map (
            O => \N__27766\,
            I => \N__27760\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27757\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__27760\,
            I => \N__27754\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__27757\,
            I => \N__27751\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27748\
        );

    \I__4427\ : Span12Mux_h
    port map (
            O => \N__27751\,
            I => \N__27745\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27742\
        );

    \I__4425\ : Span12Mux_v
    port map (
            O => \N__27745\,
            I => \N__27739\
        );

    \I__4424\ : Span12Mux_s11_v
    port map (
            O => \N__27742\,
            I => \N__27736\
        );

    \I__4423\ : Odrv12
    port map (
            O => \N__27739\,
            I => \data_index_9_N_216_7\
        );

    \I__4422\ : Odrv12
    port map (
            O => \N__27736\,
            I => \data_index_9_N_216_7\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__27731\,
            I => \n20663_cascade_\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27728\,
            I => \bfn_10_14_0_\
        );

    \I__4419\ : InMux
    port map (
            O => \N__27725\,
            I => n19384
        );

    \I__4418\ : InMux
    port map (
            O => \N__27722\,
            I => n19385
        );

    \I__4417\ : InMux
    port map (
            O => \N__27719\,
            I => n19386
        );

    \I__4416\ : InMux
    port map (
            O => \N__27716\,
            I => n19387
        );

    \I__4415\ : IoInMux
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__4413\ : Span4Mux_s2_v
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__4412\ : Sp12to4
    port map (
            O => \N__27704\,
            I => \N__27700\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27697\
        );

    \I__4410\ : Span12Mux_h
    port map (
            O => \N__27700\,
            I => \N__27694\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27690\
        );

    \I__4408\ : Span12Mux_v
    port map (
            O => \N__27694\,
            I => \N__27687\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27684\
        );

    \I__4406\ : Span4Mux_h
    port map (
            O => \N__27690\,
            I => \N__27681\
        );

    \I__4405\ : Odrv12
    port map (
            O => \N__27687\,
            I => \IAC_OSR1\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27684\,
            I => \IAC_OSR1\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__27681\,
            I => \IAC_OSR1\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27669\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27666\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27663\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__27669\,
            I => comm_cmd_4
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27666\,
            I => comm_cmd_4
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__27663\,
            I => comm_cmd_4
        );

    \I__4396\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27652\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__27655\,
            I => \N__27649\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27645\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27642\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27639\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__27645\,
            I => \N__27636\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27633\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27639\,
            I => buf_dds1_3
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__27636\,
            I => buf_dds1_3
        );

    \I__4387\ : Odrv12
    port map (
            O => \N__27633\,
            I => buf_dds1_3
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27619\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__27622\,
            I => \N__27616\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__27619\,
            I => \N__27612\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27609\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27615\,
            I => \N__27606\
        );

    \I__4380\ : Span4Mux_h
    port map (
            O => \N__27612\,
            I => \N__27603\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__27609\,
            I => \N__27600\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27606\,
            I => \N__27597\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__27603\,
            I => \N__27592\
        );

    \I__4376\ : Span4Mux_v
    port map (
            O => \N__27600\,
            I => \N__27587\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__27597\,
            I => \N__27587\
        );

    \I__4374\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27584\
        );

    \I__4373\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27581\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__27592\,
            I => \buf_cfgRTD_1\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__27587\,
            I => \buf_cfgRTD_1\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__27584\,
            I => \buf_cfgRTD_1\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27581\,
            I => \buf_cfgRTD_1\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27566\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27566\,
            I => \N__27563\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__27563\,
            I => \N__27559\
        );

    \I__4364\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27556\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__27559\,
            I => \buf_readRTD_9\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__27556\,
            I => \buf_readRTD_9\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__27542\,
            I => n9_adj_1416
        );

    \I__4357\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27534\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27531\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__27537\,
            I => \N__27528\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27534\,
            I => \N__27525\
        );

    \I__4353\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27522\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27519\
        );

    \I__4351\ : Span12Mux_v
    port map (
            O => \N__27525\,
            I => \N__27516\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27513\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__27519\,
            I => buf_dds1_0
        );

    \I__4348\ : Odrv12
    port map (
            O => \N__27516\,
            I => buf_dds1_0
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__27513\,
            I => buf_dds1_0
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__27506\,
            I => \N__27502\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__27505\,
            I => \N__27498\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27495\
        );

    \I__4343\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27492\
        );

    \I__4342\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27489\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27484\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27492\,
            I => \N__27484\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27489\,
            I => \N__27480\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__27484\,
            I => \N__27477\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \N__27474\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__27480\,
            I => \N__27468\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__27477\,
            I => \N__27468\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27465\
        );

    \I__4333\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27462\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__27468\,
            I => \buf_cfgRTD_5\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27465\,
            I => \buf_cfgRTD_5\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27462\,
            I => \buf_cfgRTD_5\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__27452\,
            I => \N__27448\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27444\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__27448\,
            I => \N__27441\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__27447\,
            I => \N__27438\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27435\
        );

    \I__4323\ : Sp12to4
    port map (
            O => \N__27441\,
            I => \N__27432\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27429\
        );

    \I__4321\ : Span4Mux_h
    port map (
            O => \N__27435\,
            I => \N__27426\
        );

    \I__4320\ : Span12Mux_h
    port map (
            O => \N__27432\,
            I => \N__27423\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__27429\,
            I => buf_adcdata_iac_18
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__27426\,
            I => buf_adcdata_iac_18
        );

    \I__4317\ : Odrv12
    port map (
            O => \N__27423\,
            I => buf_adcdata_iac_18
        );

    \I__4316\ : IoInMux
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__27413\,
            I => \N__27410\
        );

    \I__4314\ : IoSpan4Mux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4313\ : Span4Mux_s2_v
    port map (
            O => \N__27407\,
            I => \N__27404\
        );

    \I__4312\ : Sp12to4
    port map (
            O => \N__27404\,
            I => \N__27400\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27396\
        );

    \I__4310\ : Span12Mux_v
    port map (
            O => \N__27400\,
            I => \N__27393\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27390\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27387\
        );

    \I__4307\ : Odrv12
    port map (
            O => \N__27393\,
            I => \IAC_FLT0\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__27390\,
            I => \IAC_FLT0\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__27387\,
            I => \IAC_FLT0\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27380\,
            I => \N__27377\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__27377\,
            I => n20825
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__27374\,
            I => \N__27371\
        );

    \I__4301\ : CascadeBuf
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__4299\ : CascadeBuf
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__4297\ : CascadeBuf
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4295\ : CascadeBuf
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4293\ : CascadeBuf
    port map (
            O => \N__27347\,
            I => \N__27344\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4291\ : CascadeBuf
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__27338\,
            I => \N__27335\
        );

    \I__4289\ : CascadeBuf
    port map (
            O => \N__27335\,
            I => \N__27332\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4287\ : CascadeBuf
    port map (
            O => \N__27329\,
            I => \N__27325\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__27328\,
            I => \N__27322\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__27325\,
            I => \N__27319\
        );

    \I__4284\ : CascadeBuf
    port map (
            O => \N__27322\,
            I => \N__27316\
        );

    \I__4283\ : CascadeBuf
    port map (
            O => \N__27319\,
            I => \N__27313\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__27316\,
            I => \N__27310\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__27313\,
            I => \N__27307\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27304\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27301\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27298\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27301\,
            I => \N__27295\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__27298\,
            I => \N__27292\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__27295\,
            I => \N__27289\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__27292\,
            I => \N__27286\
        );

    \I__4273\ : Sp12to4
    port map (
            O => \N__27289\,
            I => \N__27283\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__27286\,
            I => \N__27280\
        );

    \I__4271\ : Span12Mux_h
    port map (
            O => \N__27283\,
            I => \N__27277\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__27280\,
            I => \data_index_9_N_216_0\
        );

    \I__4269\ : Odrv12
    port map (
            O => \N__27277\,
            I => \data_index_9_N_216_0\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27265\
        );

    \I__4267\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27265\
        );

    \I__4266\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27262\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__27265\,
            I => comm_cmd_5
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__27262\,
            I => comm_cmd_5
        );

    \I__4263\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27252\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27249\
        );

    \I__4261\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27246\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27252\,
            I => comm_cmd_6
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__27249\,
            I => comm_cmd_6
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__27246\,
            I => comm_cmd_6
        );

    \I__4257\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__27233\,
            I => \N__27229\
        );

    \I__4254\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27226\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__27229\,
            I => cmd_rdadcbuf_31
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__27226\,
            I => cmd_rdadcbuf_31
        );

    \I__4251\ : InMux
    port map (
            O => \N__27221\,
            I => \ADC_VDC.n19452\
        );

    \I__4250\ : CascadeMux
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__4249\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__27209\,
            I => \N__27205\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__27205\,
            I => cmd_rdadcbuf_32
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__27202\,
            I => cmd_rdadcbuf_32
        );

    \I__4243\ : InMux
    port map (
            O => \N__27197\,
            I => \bfn_10_9_0_\
        );

    \I__4242\ : InMux
    port map (
            O => \N__27194\,
            I => \ADC_VDC.n19454\
        );

    \I__4241\ : CEMux
    port map (
            O => \N__27191\,
            I => \N__27187\
        );

    \I__4240\ : CEMux
    port map (
            O => \N__27190\,
            I => \N__27184\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__27187\,
            I => \N__27180\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__27184\,
            I => \N__27177\
        );

    \I__4237\ : CEMux
    port map (
            O => \N__27183\,
            I => \N__27174\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__27180\,
            I => \N__27166\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__27177\,
            I => \N__27166\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27163\
        );

    \I__4233\ : CEMux
    port map (
            O => \N__27173\,
            I => \N__27160\
        );

    \I__4232\ : CEMux
    port map (
            O => \N__27172\,
            I => \N__27156\
        );

    \I__4231\ : CEMux
    port map (
            O => \N__27171\,
            I => \N__27153\
        );

    \I__4230\ : Span4Mux_h
    port map (
            O => \N__27166\,
            I => \N__27148\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__27163\,
            I => \N__27148\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27145\
        );

    \I__4227\ : CEMux
    port map (
            O => \N__27159\,
            I => \N__27142\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27156\,
            I => \N__27139\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__27153\,
            I => \N__27136\
        );

    \I__4224\ : Span4Mux_h
    port map (
            O => \N__27148\,
            I => \N__27133\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__27145\,
            I => \N__27130\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27142\,
            I => \N__27127\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__27139\,
            I => \N__27124\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__27136\,
            I => \N__27117\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__27133\,
            I => \N__27117\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__27130\,
            I => \N__27117\
        );

    \I__4217\ : Span4Mux_h
    port map (
            O => \N__27127\,
            I => \N__27114\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__27124\,
            I => \ADC_VDC.n13038\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__27117\,
            I => \ADC_VDC.n13038\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__27114\,
            I => \ADC_VDC.n13038\
        );

    \I__4213\ : SRMux
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__4212\ : SRMux
    port map (
            O => \N__27106\,
            I => \N__27096\
        );

    \I__4211\ : SRMux
    port map (
            O => \N__27105\,
            I => \N__27092\
        );

    \I__4210\ : SRMux
    port map (
            O => \N__27104\,
            I => \N__27089\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27101\,
            I => \N__27086\
        );

    \I__4208\ : SRMux
    port map (
            O => \N__27100\,
            I => \N__27083\
        );

    \I__4207\ : SRMux
    port map (
            O => \N__27099\,
            I => \N__27080\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27096\,
            I => \N__27077\
        );

    \I__4205\ : SRMux
    port map (
            O => \N__27095\,
            I => \N__27074\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27071\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__27089\,
            I => \N__27066\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__27086\,
            I => \N__27066\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27063\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__27080\,
            I => \N__27060\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__27077\,
            I => \N__27055\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27055\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__27071\,
            I => \N__27052\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__27066\,
            I => \N__27047\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__27063\,
            I => \N__27047\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__27060\,
            I => \N__27044\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__27055\,
            I => \N__27041\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__27052\,
            I => \N__27038\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__27047\,
            I => \ADC_VDC.n14931\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__27044\,
            I => \ADC_VDC.n14931\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__27041\,
            I => \ADC_VDC.n14931\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__27038\,
            I => \ADC_VDC.n14931\
        );

    \I__4187\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__4185\ : Span12Mux_h
    port map (
            O => \N__27023\,
            I => \N__27018\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27015\
        );

    \I__4183\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27012\
        );

    \I__4182\ : Odrv12
    port map (
            O => \N__27018\,
            I => cmd_rdadcbuf_34
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__27015\,
            I => cmd_rdadcbuf_34
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__27012\,
            I => cmd_rdadcbuf_34
        );

    \I__4179\ : InMux
    port map (
            O => \N__27005\,
            I => \ADC_VDC.n19455\
        );

    \I__4178\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26999\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__26999\,
            I => \ADC_VDC.cmd_rdadcbuf_35_N_1139_34\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__4175\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26987\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__26987\,
            I => \N__26984\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__26981\,
            I => n20824
        );

    \I__4170\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26975\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__26975\,
            I => n22118
        );

    \I__4168\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26967\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__26971\,
            I => \N__26964\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26961\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26958\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26955\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26961\,
            I => cmd_rdadctmp_8
        );

    \I__4162\ : Odrv12
    port map (
            O => \N__26958\,
            I => cmd_rdadctmp_8
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26955\,
            I => cmd_rdadctmp_8
        );

    \I__4160\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26944\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26941\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__26944\,
            I => cmd_rdadcbuf_22
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26941\,
            I => cmd_rdadcbuf_22
        );

    \I__4156\ : InMux
    port map (
            O => \N__26936\,
            I => \ADC_VDC.n19443\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26930\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__26930\,
            I => \N__26926\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26923\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__26926\,
            I => cmd_rdadcbuf_23
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26923\,
            I => cmd_rdadcbuf_23
        );

    \I__4150\ : InMux
    port map (
            O => \N__26918\,
            I => \ADC_VDC.n19444\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26915\,
            I => \bfn_10_8_0_\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26912\,
            I => \ADC_VDC.n19446\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26909\,
            I => \ADC_VDC.n19447\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26906\,
            I => \ADC_VDC.n19448\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26897\,
            I => \N__26894\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__26894\,
            I => \N__26890\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26887\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__26890\,
            I => cmd_rdadcbuf_28
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26887\,
            I => cmd_rdadcbuf_28
        );

    \I__4138\ : InMux
    port map (
            O => \N__26882\,
            I => \ADC_VDC.n19449\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26872\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26869\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__26872\,
            I => cmd_rdadcbuf_29
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26869\,
            I => cmd_rdadcbuf_29
        );

    \I__4132\ : InMux
    port map (
            O => \N__26864\,
            I => \ADC_VDC.n19450\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26854\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26851\
        );

    \I__4128\ : Odrv12
    port map (
            O => \N__26854\,
            I => cmd_rdadcbuf_30
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26851\,
            I => cmd_rdadcbuf_30
        );

    \I__4126\ : InMux
    port map (
            O => \N__26846\,
            I => \ADC_VDC.n19451\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26838\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26835\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26832\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26838\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26835\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26832\,
            I => cmd_rdadctmp_14_adj_1465
        );

    \I__4119\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26821\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__26824\,
            I => \N__26818\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26821\,
            I => \N__26815\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26812\
        );

    \I__4115\ : Odrv12
    port map (
            O => \N__26815\,
            I => cmd_rdadcbuf_14
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__26812\,
            I => cmd_rdadcbuf_14
        );

    \I__4113\ : InMux
    port map (
            O => \N__26807\,
            I => \ADC_VDC.n19435\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__26804\,
            I => \N__26799\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26794\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26794\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26791\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26794\,
            I => cmd_rdadctmp_15_adj_1464
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26791\,
            I => cmd_rdadctmp_15_adj_1464
        );

    \I__4106\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26779\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26776\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__26779\,
            I => cmd_rdadcbuf_15
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26776\,
            I => cmd_rdadcbuf_15
        );

    \I__4101\ : InMux
    port map (
            O => \N__26771\,
            I => \ADC_VDC.n19436\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__26768\,
            I => \N__26763\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__26767\,
            I => \N__26760\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__26766\,
            I => \N__26757\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26752\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26752\
        );

    \I__4095\ : InMux
    port map (
            O => \N__26757\,
            I => \N__26749\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26752\,
            I => cmd_rdadctmp_16_adj_1463
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26749\,
            I => cmd_rdadctmp_16_adj_1463
        );

    \I__4092\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__26738\,
            I => \N__26734\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26731\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__26734\,
            I => cmd_rdadcbuf_16
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26731\,
            I => cmd_rdadcbuf_16
        );

    \I__4086\ : InMux
    port map (
            O => \N__26726\,
            I => \bfn_10_7_0_\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__26723\,
            I => \N__26718\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26713\
        );

    \I__4083\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26713\
        );

    \I__4082\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26710\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__26713\,
            I => cmd_rdadctmp_17_adj_1462
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__26710\,
            I => cmd_rdadctmp_17_adj_1462
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__26705\,
            I => \N__26702\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__26696\,
            I => \N__26692\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26689\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__26692\,
            I => cmd_rdadcbuf_17
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26689\,
            I => cmd_rdadcbuf_17
        );

    \I__4072\ : InMux
    port map (
            O => \N__26684\,
            I => \ADC_VDC.n19438\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__26681\,
            I => \N__26676\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26673\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26670\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26667\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26673\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26670\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__26667\,
            I => cmd_rdadctmp_18_adj_1461
        );

    \I__4064\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__26654\,
            I => \N__26650\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26647\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26650\,
            I => cmd_rdadcbuf_18
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__26647\,
            I => cmd_rdadcbuf_18
        );

    \I__4058\ : InMux
    port map (
            O => \N__26642\,
            I => \ADC_VDC.n19439\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26634\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26629\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26629\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26626\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26629\,
            I => cmd_rdadctmp_19_adj_1460
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26626\,
            I => cmd_rdadctmp_19_adj_1460
        );

    \I__4051\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__26618\,
            I => \N__26614\
        );

    \I__4049\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__4048\ : Odrv12
    port map (
            O => \N__26614\,
            I => cmd_rdadcbuf_19
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__26611\,
            I => cmd_rdadcbuf_19
        );

    \I__4046\ : InMux
    port map (
            O => \N__26606\,
            I => \ADC_VDC.n19440\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__26603\,
            I => \N__26598\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26595\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26592\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26589\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26586\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26583\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__26589\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__26586\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26583\,
            I => cmd_rdadctmp_20_adj_1459
        );

    \I__4036\ : InMux
    port map (
            O => \N__26576\,
            I => \ADC_VDC.n19441\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__26573\,
            I => \N__26570\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26565\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26560\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26560\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26557\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__26560\,
            I => cmd_rdadctmp_21_adj_1458
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__26557\,
            I => cmd_rdadctmp_21_adj_1458
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__26543\,
            I => \N__26539\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26536\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__26539\,
            I => cmd_rdadcbuf_21
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__26536\,
            I => cmd_rdadcbuf_21
        );

    \I__4021\ : InMux
    port map (
            O => \N__26531\,
            I => \ADC_VDC.n19442\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26528\,
            I => \ADC_VDC.n19427\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26521\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \N__26517\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__26521\,
            I => \N__26514\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26520\,
            I => \N__26511\
        );

    \I__4015\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26508\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__26514\,
            I => cmd_rdadctmp_7_adj_1472
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__26511\,
            I => cmd_rdadctmp_7_adj_1472
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__26508\,
            I => cmd_rdadctmp_7_adj_1472
        );

    \I__4011\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__26498\,
            I => \ADC_VDC.cmd_rdadcbuf_7\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26495\,
            I => \ADC_VDC.n19428\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26488\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__26491\,
            I => \N__26484\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26488\,
            I => \N__26481\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26478\
        );

    \I__4004\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26475\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__26481\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__26478\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__26475\,
            I => cmd_rdadctmp_8_adj_1471
        );

    \I__4000\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__26465\,
            I => \ADC_VDC.cmd_rdadcbuf_8\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26462\,
            I => \bfn_10_6_0_\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \N__26455\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__26458\,
            I => \N__26451\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26448\
        );

    \I__3994\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26445\
        );

    \I__3993\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26442\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__26448\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__26445\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26442\,
            I => cmd_rdadctmp_9_adj_1470
        );

    \I__3989\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__26432\,
            I => \ADC_VDC.cmd_rdadcbuf_9\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26429\,
            I => \ADC_VDC.n19430\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__26426\,
            I => \N__26422\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__26425\,
            I => \N__26418\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26415\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26412\
        );

    \I__3982\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26409\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__26415\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__26412\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26409\,
            I => cmd_rdadctmp_10_adj_1469
        );

    \I__3978\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__26399\,
            I => \ADC_VDC.cmd_rdadcbuf_10\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26396\,
            I => \ADC_VDC.n19431\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__26393\,
            I => \N__26388\
        );

    \I__3974\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26383\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26383\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26380\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26383\,
            I => cmd_rdadctmp_11_adj_1468
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__26380\,
            I => cmd_rdadctmp_11_adj_1468
        );

    \I__3969\ : InMux
    port map (
            O => \N__26375\,
            I => \ADC_VDC.n19432\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26368\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__26371\,
            I => \N__26365\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26361\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26356\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26356\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26353\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26356\,
            I => cmd_rdadctmp_12_adj_1467
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__26353\,
            I => cmd_rdadctmp_12_adj_1467
        );

    \I__3960\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__26345\,
            I => \N__26341\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26338\
        );

    \I__3957\ : Odrv12
    port map (
            O => \N__26341\,
            I => cmd_rdadcbuf_12
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__26338\,
            I => cmd_rdadcbuf_12
        );

    \I__3955\ : InMux
    port map (
            O => \N__26333\,
            I => \ADC_VDC.n19433\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26323\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26323\
        );

    \I__3952\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26320\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26323\,
            I => cmd_rdadctmp_13_adj_1466
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26320\,
            I => cmd_rdadctmp_13_adj_1466
        );

    \I__3949\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26308\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \N__26305\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__26308\,
            I => \N__26302\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26299\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__26302\,
            I => cmd_rdadcbuf_13
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__26299\,
            I => cmd_rdadcbuf_13
        );

    \I__3942\ : InMux
    port map (
            O => \N__26294\,
            I => \ADC_VDC.n19434\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__26291\,
            I => \N__26285\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__26290\,
            I => \N__26281\
        );

    \I__3939\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26262\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26262\
        );

    \I__3937\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26262\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26262\
        );

    \I__3935\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26262\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__26280\,
            I => \N__26259\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__26279\,
            I => \N__26256\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__26278\,
            I => \N__26251\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__26277\,
            I => \N__26247\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__26276\,
            I => \N__26243\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__26275\,
            I => \N__26237\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__26274\,
            I => \N__26233\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__26273\,
            I => \N__26229\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26226\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26215\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26215\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26215\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26215\
        );

    \I__3921\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26215\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26202\
        );

    \I__3919\ : InMux
    port map (
            O => \N__26247\,
            I => \N__26202\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26202\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26202\
        );

    \I__3916\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26202\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26202\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26189\
        );

    \I__3913\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26189\
        );

    \I__3912\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26189\
        );

    \I__3911\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26189\
        );

    \I__3910\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26189\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26189\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__26226\,
            I => n12875
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__26215\,
            I => n12875
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26202\,
            I => n12875
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__26189\,
            I => n12875
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26176\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__26179\,
            I => \N__26172\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26167\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26167\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26164\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__26167\,
            I => cmd_rdadctmp_0_adj_1479
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__26164\,
            I => cmd_rdadctmp_0_adj_1479
        );

    \I__3897\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__26156\,
            I => \ADC_VDC.cmd_rdadcbuf_0\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__26153\,
            I => \N__26148\
        );

    \I__3894\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26145\
        );

    \I__3893\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26142\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26139\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__26145\,
            I => cmd_rdadctmp_1_adj_1478
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__26142\,
            I => cmd_rdadctmp_1_adj_1478
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__26139\,
            I => cmd_rdadctmp_1_adj_1478
        );

    \I__3888\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26129\,
            I => \ADC_VDC.cmd_rdadcbuf_1\
        );

    \I__3886\ : InMux
    port map (
            O => \N__26126\,
            I => \ADC_VDC.n19422\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__26123\,
            I => \N__26118\
        );

    \I__3884\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26113\
        );

    \I__3883\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26113\
        );

    \I__3882\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26110\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__26113\,
            I => cmd_rdadctmp_2_adj_1477
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__26110\,
            I => cmd_rdadctmp_2_adj_1477
        );

    \I__3879\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__26102\,
            I => \ADC_VDC.cmd_rdadcbuf_2\
        );

    \I__3877\ : InMux
    port map (
            O => \N__26099\,
            I => \ADC_VDC.n19423\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__26096\,
            I => \N__26092\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__26095\,
            I => \N__26088\
        );

    \I__3874\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26083\
        );

    \I__3873\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26083\
        );

    \I__3872\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26080\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__26083\,
            I => cmd_rdadctmp_3_adj_1476
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__26080\,
            I => cmd_rdadctmp_3_adj_1476
        );

    \I__3869\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__26072\,
            I => \ADC_VDC.cmd_rdadcbuf_3\
        );

    \I__3867\ : InMux
    port map (
            O => \N__26069\,
            I => \ADC_VDC.n19424\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__26066\,
            I => \N__26061\
        );

    \I__3865\ : InMux
    port map (
            O => \N__26065\,
            I => \N__26058\
        );

    \I__3864\ : InMux
    port map (
            O => \N__26064\,
            I => \N__26055\
        );

    \I__3863\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26052\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__26058\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__26055\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__26052\,
            I => cmd_rdadctmp_4_adj_1475
        );

    \I__3859\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__26042\,
            I => \ADC_VDC.cmd_rdadcbuf_4\
        );

    \I__3857\ : InMux
    port map (
            O => \N__26039\,
            I => \ADC_VDC.n19425\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__26036\,
            I => \N__26032\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__26035\,
            I => \N__26028\
        );

    \I__3854\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26025\
        );

    \I__3853\ : InMux
    port map (
            O => \N__26031\,
            I => \N__26022\
        );

    \I__3852\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26019\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__26025\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__26022\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__26019\,
            I => cmd_rdadctmp_5_adj_1474
        );

    \I__3848\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__26009\,
            I => \ADC_VDC.cmd_rdadcbuf_5\
        );

    \I__3846\ : InMux
    port map (
            O => \N__26006\,
            I => \ADC_VDC.n19426\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \N__25998\
        );

    \I__3844\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25993\
        );

    \I__3843\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25993\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25990\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__25993\,
            I => cmd_rdadctmp_6_adj_1473
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25990\,
            I => cmd_rdadctmp_6_adj_1473
        );

    \I__3839\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25982\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25982\,
            I => \ADC_VDC.cmd_rdadcbuf_6\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25973\,
            I => \N__25969\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25965\
        );

    \I__3833\ : Span4Mux_h
    port map (
            O => \N__25969\,
            I => \N__25962\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25959\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25965\,
            I => cmd_rdadctmp_12
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__25962\,
            I => cmd_rdadctmp_12
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25959\,
            I => cmd_rdadctmp_12
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25945\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__25948\,
            I => \N__25941\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__25945\,
            I => \N__25938\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25935\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25932\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__25938\,
            I => \N__25927\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25927\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__25932\,
            I => cmd_rdadctmp_13
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__25927\,
            I => cmd_rdadctmp_13
        );

    \I__3818\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25918\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25918\,
            I => \N__25912\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25909\
        );

    \I__3814\ : Span4Mux_h
    port map (
            O => \N__25912\,
            I => \N__25906\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25909\,
            I => cmd_rdadctmp_6
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__25906\,
            I => cmd_rdadctmp_6
        );

    \I__3811\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25897\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25897\,
            I => cmd_rdadctmp_7
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25894\,
            I => cmd_rdadctmp_7
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25882\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__25885\,
            I => \N__25879\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25882\,
            I => \N__25875\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25870\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25878\,
            I => \N__25870\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__25875\,
            I => cmd_rdadctmp_13_adj_1437
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25870\,
            I => cmd_rdadctmp_13_adj_1437
        );

    \I__3799\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25857\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25854\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25851\
        );

    \I__3795\ : Span4Mux_h
    port map (
            O => \N__25857\,
            I => \N__25846\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25846\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25851\,
            I => buf_adcdata_iac_5
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__25846\,
            I => buf_adcdata_iac_5
        );

    \I__3791\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__25832\,
            I => buf_data_iac_5
        );

    \I__3787\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25826\,
            I => \N__25823\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__25823\,
            I => n22_adj_1632
        );

    \I__3784\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25817\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__3781\ : Span4Mux_h
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__25808\,
            I => \ADC_VDC.n21718\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__25805\,
            I => \n12383_cascade_\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25794\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25791\
        );

    \I__3775\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25788\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__25794\,
            I => buf_dds1_10
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__25791\,
            I => buf_dds1_10
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25788\,
            I => buf_dds1_10
        );

    \I__3771\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25777\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25774\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25777\,
            I => n20673
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25774\,
            I => n20673
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__25769\,
            I => \n11412_cascade_\
        );

    \I__3766\ : IoInMux
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__3764\ : IoSpan4Mux
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__3763\ : IoSpan4Mux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__3762\ : Span4Mux_s2_v
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__25748\,
            I => \AC_ADC_SYNC\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25741\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25737\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__25741\,
            I => \N__25734\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25731\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25737\,
            I => buf_dds1_4
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__25734\,
            I => buf_dds1_4
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__25731\,
            I => buf_dds1_4
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__25724\,
            I => \n8_adj_1555_cascade_\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__3750\ : CascadeBuf
    port map (
            O => \N__25718\,
            I => \N__25715\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \N__25712\
        );

    \I__3748\ : CascadeBuf
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__3746\ : CascadeBuf
    port map (
            O => \N__25706\,
            I => \N__25703\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__3744\ : CascadeBuf
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3742\ : CascadeBuf
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__3740\ : CascadeBuf
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__3738\ : CascadeBuf
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__3736\ : CascadeBuf
    port map (
            O => \N__25676\,
            I => \N__25672\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__25675\,
            I => \N__25669\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25666\
        );

    \I__3733\ : CascadeBuf
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__3732\ : CascadeBuf
    port map (
            O => \N__25666\,
            I => \N__25660\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__25663\,
            I => \N__25657\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25651\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25648\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__3725\ : Span12Mux_h
    port map (
            O => \N__25645\,
            I => \N__25639\
        );

    \I__3724\ : Span12Mux_v
    port map (
            O => \N__25642\,
            I => \N__25636\
        );

    \I__3723\ : Span12Mux_v
    port map (
            O => \N__25639\,
            I => \N__25633\
        );

    \I__3722\ : Span12Mux_h
    port map (
            O => \N__25636\,
            I => \N__25630\
        );

    \I__3721\ : Odrv12
    port map (
            O => \N__25633\,
            I => \data_index_9_N_216_8\
        );

    \I__3720\ : Odrv12
    port map (
            O => \N__25630\,
            I => \data_index_9_N_216_8\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25622\,
            I => n8_adj_1555
        );

    \I__3717\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25616\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__25613\,
            I => n22040
        );

    \I__3714\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25605\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25602\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25599\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__25605\,
            I => buf_dds1_9
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__25602\,
            I => buf_dds1_9
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__25599\,
            I => buf_dds1_9
        );

    \I__3708\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25588\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25584\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25588\,
            I => \N__25581\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25578\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25584\,
            I => buf_dds1_8
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__25581\,
            I => buf_dds1_8
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25578\,
            I => buf_dds1_8
        );

    \I__3701\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__25568\,
            I => n20849
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__3698\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25559\,
            I => n22103
        );

    \I__3696\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__3693\ : Sp12to4
    port map (
            O => \N__25547\,
            I => \N__25542\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \N__25539\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25536\
        );

    \I__3690\ : Span12Mux_h
    port map (
            O => \N__25542\,
            I => \N__25533\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25530\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25536\,
            I => buf_adcdata_iac_17
        );

    \I__3687\ : Odrv12
    port map (
            O => \N__25533\,
            I => buf_adcdata_iac_17
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__25530\,
            I => buf_adcdata_iac_17
        );

    \I__3685\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__3683\ : Span12Mux_v
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3682\ : Span12Mux_h
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__3681\ : Odrv12
    port map (
            O => \N__25511\,
            I => buf_data_iac_21
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__25508\,
            I => \n20876_cascade_\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25502\,
            I => n22106
        );

    \I__3677\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__25496\,
            I => n20875
        );

    \I__3675\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25490\,
            I => n22022
        );

    \I__3673\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25484\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25480\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25477\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__25480\,
            I => \N__25474\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25477\,
            I => \N__25471\
        );

    \I__3668\ : Sp12to4
    port map (
            O => \N__25474\,
            I => \N__25467\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__25471\,
            I => \N__25464\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25470\,
            I => \N__25461\
        );

    \I__3665\ : Span12Mux_h
    port map (
            O => \N__25467\,
            I => \N__25458\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__25464\,
            I => \N__25455\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__25461\,
            I => buf_adcdata_vac_21
        );

    \I__3662\ : Odrv12
    port map (
            O => \N__25458\,
            I => buf_adcdata_vac_21
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__25455\,
            I => buf_adcdata_vac_21
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__25448\,
            I => \N__25445\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__25439\,
            I => \N__25436\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__25436\,
            I => \N__25432\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25429\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__25432\,
            I => buf_adcdata_vdc_21
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25429\,
            I => buf_adcdata_vdc_21
        );

    \I__3652\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__25421\,
            I => n22184
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__25409\,
            I => \N__25405\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25402\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__25405\,
            I => \buf_readRTD_12\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__25402\,
            I => \buf_readRTD_12\
        );

    \I__3643\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__25388\,
            I => n22202
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__25376\,
            I => \N__25372\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25369\
        );

    \I__3634\ : Odrv4
    port map (
            O => \N__25372\,
            I => \buf_readRTD_8\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25369\,
            I => \buf_readRTD_8\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__25364\,
            I => \N__25361\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25356\
        );

    \I__3630\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25353\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \N__25350\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25347\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__25353\,
            I => \N__25344\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25341\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__25347\,
            I => \N__25333\
        );

    \I__3624\ : Span4Mux_h
    port map (
            O => \N__25344\,
            I => \N__25333\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25333\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25329\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__25333\,
            I => \N__25326\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25323\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25329\,
            I => \N__25320\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__25326\,
            I => \buf_cfgRTD_0\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__25323\,
            I => \buf_cfgRTD_0\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__25320\,
            I => \buf_cfgRTD_0\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__25298\,
            I => \N__25293\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25290\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25287\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__25293\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25290\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__25287\,
            I => cmd_rdadctmp_27_adj_1423
        );

    \I__3604\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25277\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__25277\,
            I => \N__25272\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25269\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25266\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__25272\,
            I => \N__25261\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25261\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25266\,
            I => buf_dds1_15
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__25261\,
            I => buf_dds1_15
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__25256\,
            I => \N__25252\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25245\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25242\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__25248\,
            I => \N__25239\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25236\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__25242\,
            I => \N__25233\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25230\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__25236\,
            I => \N__25225\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__25233\,
            I => \N__25220\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25230\,
            I => \N__25220\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25217\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25214\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__25225\,
            I => \buf_cfgRTD_4\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__25220\,
            I => \buf_cfgRTD_4\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__25217\,
            I => \buf_cfgRTD_4\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25214\,
            I => \buf_cfgRTD_4\
        );

    \I__3579\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25201\
        );

    \I__3578\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25198\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25191\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__25198\,
            I => \N__25191\
        );

    \I__3575\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25188\
        );

    \I__3574\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25184\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__25191\,
            I => \N__25181\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25188\,
            I => \N__25178\
        );

    \I__3571\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25175\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__25184\,
            I => \N__25172\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__25181\,
            I => \buf_cfgRTD_3\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__25178\,
            I => \buf_cfgRTD_3\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25175\,
            I => \buf_cfgRTD_3\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__25172\,
            I => \buf_cfgRTD_3\
        );

    \I__3565\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25160\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25156\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__25159\,
            I => \N__25153\
        );

    \I__3562\ : Span4Mux_h
    port map (
            O => \N__25156\,
            I => \N__25150\
        );

    \I__3561\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25147\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__25150\,
            I => cmd_rdadctmp_7_adj_1443
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__25147\,
            I => cmd_rdadctmp_7_adj_1443
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__3557\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__25133\,
            I => \N__25129\
        );

    \I__3554\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__25129\,
            I => \buf_readRTD_13\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__25126\,
            I => \buf_readRTD_13\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25117\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25114\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25117\,
            I => \N__25111\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__25114\,
            I => \N__25108\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__25111\,
            I => \buf_readRTD_10\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__25108\,
            I => \buf_readRTD_10\
        );

    \I__3545\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25099\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__25102\,
            I => \N__25096\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25092\
        );

    \I__3542\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25089\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__25095\,
            I => \N__25086\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__25092\,
            I => \N__25081\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25078\
        );

    \I__3538\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25075\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25072\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25069\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__25081\,
            I => \buf_cfgRTD_2\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__25078\,
            I => \buf_cfgRTD_2\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__25075\,
            I => \buf_cfgRTD_2\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__25072\,
            I => \buf_cfgRTD_2\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__25069\,
            I => \buf_cfgRTD_2\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__25052\,
            I => n20834
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__25049\,
            I => \N__25044\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__25048\,
            I => \N__25041\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25035\
        );

    \I__3524\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25027\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25024\
        );

    \I__3522\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25021\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25006\
        );

    \I__3520\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25003\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__25035\,
            I => \N__25000\
        );

    \I__3518\ : InMux
    port map (
            O => \N__25034\,
            I => \N__24989\
        );

    \I__3517\ : InMux
    port map (
            O => \N__25033\,
            I => \N__24989\
        );

    \I__3516\ : InMux
    port map (
            O => \N__25032\,
            I => \N__24989\
        );

    \I__3515\ : InMux
    port map (
            O => \N__25031\,
            I => \N__24989\
        );

    \I__3514\ : InMux
    port map (
            O => \N__25030\,
            I => \N__24989\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__25027\,
            I => \N__24984\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__24984\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__24981\
        );

    \I__3510\ : InMux
    port map (
            O => \N__25020\,
            I => \N__24976\
        );

    \I__3509\ : InMux
    port map (
            O => \N__25019\,
            I => \N__24976\
        );

    \I__3508\ : InMux
    port map (
            O => \N__25018\,
            I => \N__24969\
        );

    \I__3507\ : InMux
    port map (
            O => \N__25017\,
            I => \N__24969\
        );

    \I__3506\ : InMux
    port map (
            O => \N__25016\,
            I => \N__24969\
        );

    \I__3505\ : InMux
    port map (
            O => \N__25015\,
            I => \N__24960\
        );

    \I__3504\ : InMux
    port map (
            O => \N__25014\,
            I => \N__24960\
        );

    \I__3503\ : InMux
    port map (
            O => \N__25013\,
            I => \N__24960\
        );

    \I__3502\ : InMux
    port map (
            O => \N__25012\,
            I => \N__24960\
        );

    \I__3501\ : InMux
    port map (
            O => \N__25011\,
            I => \N__24953\
        );

    \I__3500\ : InMux
    port map (
            O => \N__25010\,
            I => \N__24953\
        );

    \I__3499\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24953\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24944\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24944\
        );

    \I__3496\ : Span4Mux_h
    port map (
            O => \N__25000\,
            I => \N__24944\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24944\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__24984\,
            I => adc_state_1_adj_1483
        );

    \I__3493\ : Odrv4
    port map (
            O => \N__24981\,
            I => adc_state_1_adj_1483
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24976\,
            I => adc_state_1_adj_1483
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24969\,
            I => adc_state_1_adj_1483
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24960\,
            I => adc_state_1_adj_1483
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24953\,
            I => adc_state_1_adj_1483
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__24944\,
            I => adc_state_1_adj_1483
        );

    \I__3487\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24925\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24925\,
            I => \RTD.n20656\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24922\,
            I => \RTD.n20656\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__24917\,
            I => \n12397_cascade_\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24908\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__24908\,
            I => \RTD.n10\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24901\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24901\,
            I => \RTD.cfg_buf_2\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24898\,
            I => \RTD.cfg_buf_2\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24889\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24886\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24889\,
            I => \N__24882\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24886\,
            I => \N__24879\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24876\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__24882\,
            I => \N__24871\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__24879\,
            I => \N__24871\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24876\,
            I => read_buf_0
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__24871\,
            I => read_buf_0
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__24866\,
            I => \N__24860\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__24865\,
            I => \N__24857\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24854\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__24863\,
            I => \N__24851\
        );

    \I__3462\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24826\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24826\
        );

    \I__3460\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24826\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24851\,
            I => \N__24826\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24826\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24826\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24823\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24814\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24814\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24814\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24814\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24809\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24809\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24786\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24786\
        );

    \I__3447\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24786\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24781\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__24823\,
            I => \N__24781\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24814\,
            I => \N__24776\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24776\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24773\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__24807\,
            I => \N__24770\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__24806\,
            I => \N__24766\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24756\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24756\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24756\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24756\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24751\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24751\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24748\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24745\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24742\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24739\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24736\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24731\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24731\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24724\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__24781\,
            I => \N__24724\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__24776\,
            I => \N__24724\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24721\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24716\
        );

    \I__3421\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24716\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24711\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24711\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24708\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__24751\,
            I => \RTD.adc_state_0\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24748\,
            I => \RTD.adc_state_0\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24745\,
            I => \RTD.adc_state_0\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24742\,
            I => \RTD.adc_state_0\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24739\,
            I => \RTD.adc_state_0\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24736\,
            I => \RTD.adc_state_0\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__24731\,
            I => \RTD.adc_state_0\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__24724\,
            I => \RTD.adc_state_0\
        );

    \I__3409\ : Odrv4
    port map (
            O => \N__24721\,
            I => \RTD.adc_state_0\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__24716\,
            I => \RTD.adc_state_0\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24711\,
            I => \RTD.adc_state_0\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__24708\,
            I => \RTD.adc_state_0\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__24683\,
            I => \N__24670\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__24682\,
            I => \N__24667\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__24681\,
            I => \N__24661\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__24680\,
            I => \N__24655\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__24679\,
            I => \N__24652\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__24678\,
            I => \N__24649\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__24677\,
            I => \N__24645\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24640\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__24675\,
            I => \N__24637\
        );

    \I__3396\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24631\
        );

    \I__3395\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24628\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24621\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24621\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24621\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24616\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24616\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24609\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24609\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24609\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24606\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24603\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24592\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24592\
        );

    \I__3382\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24592\
        );

    \I__3381\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24592\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24592\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24588\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24585\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24579\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24579\
        );

    \I__3375\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24574\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24574\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24571\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24568\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24561\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24561\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24561\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__24606\,
            I => \N__24554\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24554\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__24592\,
            I => \N__24554\
        );

    \I__3365\ : InMux
    port map (
            O => \N__24591\,
            I => \N__24551\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24546\
        );

    \I__3363\ : Span4Mux_v
    port map (
            O => \N__24585\,
            I => \N__24546\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24543\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24579\,
            I => \N__24538\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24538\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__24571\,
            I => \N__24529\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__24568\,
            I => \N__24529\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__24561\,
            I => \N__24529\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__24554\,
            I => \N__24529\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24551\,
            I => adc_state_3_adj_1481
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__24546\,
            I => adc_state_3_adj_1481
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24543\,
            I => adc_state_3_adj_1481
        );

    \I__3352\ : Odrv12
    port map (
            O => \N__24538\,
            I => adc_state_3_adj_1481
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__24529\,
            I => adc_state_3_adj_1481
        );

    \I__3350\ : SRMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24511\
        );

    \I__3348\ : SRMux
    port map (
            O => \N__24514\,
            I => \N__24508\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__24511\,
            I => \N__24505\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__24505\,
            I => \N__24499\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__24502\,
            I => \N__24496\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__24499\,
            I => \RTD.n14717\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__24496\,
            I => \RTD.n14717\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__24488\,
            I => n16_adj_1524
        );

    \I__3339\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24481\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24481\,
            I => \RTD.cfg_buf_4\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__24478\,
            I => \RTD.cfg_buf_4\
        );

    \I__3335\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24463\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24456\
        );

    \I__3333\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24456\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24456\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24451\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24451\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__24467\,
            I => \N__24428\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24414\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24406\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24401\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24401\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24394\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24394\
        );

    \I__3322\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24394\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24383\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24383\
        );

    \I__3319\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24383\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24444\,
            I => \N__24383\
        );

    \I__3317\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24383\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24372\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24372\
        );

    \I__3314\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24372\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24372\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24372\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24362\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24362\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24362\
        );

    \I__3308\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24351\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24351\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24351\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24351\
        );

    \I__3304\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24351\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24334\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24334\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24334\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24334\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24334\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24334\
        );

    \I__3297\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24334\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24334\
        );

    \I__3295\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24329\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24329\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24326\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24323\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24316\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24316\
        );

    \I__3289\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24316\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24311\
        );

    \I__3287\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24311\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__24406\,
            I => \N__24302\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__24401\,
            I => \N__24302\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__24394\,
            I => \N__24302\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__24383\,
            I => \N__24302\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__24372\,
            I => \N__24299\
        );

    \I__3281\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24292\
        );

    \I__3280\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24292\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24292\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24287\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24287\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__24334\,
            I => adc_state_2_adj_1482
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24329\,
            I => adc_state_2_adj_1482
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__24326\,
            I => adc_state_2_adj_1482
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__24323\,
            I => adc_state_2_adj_1482
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24316\,
            I => adc_state_2_adj_1482
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24311\,
            I => adc_state_2_adj_1482
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__24302\,
            I => adc_state_2_adj_1482
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__24299\,
            I => adc_state_2_adj_1482
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__24292\,
            I => adc_state_2_adj_1482
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__24287\,
            I => adc_state_2_adj_1482
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24255\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__24259\,
            I => \N__24252\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__24258\,
            I => \N__24249\
        );

    \I__3261\ : Span4Mux_h
    port map (
            O => \N__24255\,
            I => \N__24246\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24252\,
            I => \N__24241\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24241\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__24246\,
            I => read_buf_6
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24241\,
            I => read_buf_6
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \N__24230\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24224\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24213\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24213\
        );

    \I__3252\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24208\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24208\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24203\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24203\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24194\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24194\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24194\
        );

    \I__3245\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24185\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24185\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24185\
        );

    \I__3242\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24185\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__24213\,
            I => \N__24182\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24208\,
            I => \N__24179\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__24203\,
            I => \N__24176\
        );

    \I__3238\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24173\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24170\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24167\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24164\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__24182\,
            I => \N__24161\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__24179\,
            I => \N__24156\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__24176\,
            I => \N__24156\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__24173\,
            I => n11730
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__24170\,
            I => n11730
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__24167\,
            I => n11730
        );

    \I__3228\ : Odrv12
    port map (
            O => \N__24164\,
            I => n11730
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__24161\,
            I => n11730
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__24156\,
            I => n11730
        );

    \I__3225\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24128\
        );

    \I__3224\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24128\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24128\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24128\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24128\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24122\
        );

    \I__3219\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24115\
        );

    \I__3218\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24115\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24115\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__24122\,
            I => \RTD.n13192\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__24115\,
            I => \RTD.n13192\
        );

    \I__3214\ : InMux
    port map (
            O => \N__24110\,
            I => \N__24091\
        );

    \I__3213\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24091\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24091\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24091\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24091\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24084\
        );

    \I__3208\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24084\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24084\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__24102\,
            I => \N__24081\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24078\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24075\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24072\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__24078\,
            I => \RTD.n20631\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__24075\,
            I => \RTD.n20631\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__24072\,
            I => \RTD.n20631\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24059\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24056\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24051\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24051\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24048\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24042\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24042\
        );

    \I__3192\ : Span12Mux_v
    port map (
            O => \N__24048\,
            I => \N__24039\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24036\
        );

    \I__3190\ : Span4Mux_v
    port map (
            O => \N__24042\,
            I => \N__24033\
        );

    \I__3189\ : Odrv12
    port map (
            O => \N__24039\,
            I => \buf_cfgRTD_7\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__24036\,
            I => \buf_cfgRTD_7\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__24033\,
            I => \buf_cfgRTD_7\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__24026\,
            I => \N__24023\
        );

    \I__3185\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24019\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24016\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__24019\,
            I => \RTD.cfg_buf_7\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__24016\,
            I => \RTD.cfg_buf_7\
        );

    \I__3181\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__24005\
        );

    \I__3179\ : Odrv12
    port map (
            O => \N__24005\,
            I => \ADC_VDC.n18479\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__24002\,
            I => \ADC_VDC.n21145_cascade_\
        );

    \I__3177\ : CEMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23993\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23993\,
            I => \ADC_VDC.n13050\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__23990\,
            I => \N__23987\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23984\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23981\
        );

    \I__3171\ : Span4Mux_v
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3170\ : Span4Mux_h
    port map (
            O => \N__23978\,
            I => \N__23973\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23968\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23968\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__23973\,
            I => read_buf_10
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23968\,
            I => read_buf_10
        );

    \I__3165\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__23957\,
            I => \N__23953\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__23956\,
            I => \N__23950\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__23953\,
            I => \N__23947\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23944\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__23947\,
            I => buf_adcdata_vdc_18
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23944\,
            I => buf_adcdata_vdc_18
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__23939\,
            I => \n20833_cascade_\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23930\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23927\
        );

    \I__3153\ : Span4Mux_h
    port map (
            O => \N__23927\,
            I => \N__23922\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23917\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23917\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__23922\,
            I => read_buf_14
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23917\,
            I => read_buf_14
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__23903\,
            I => \N__23899\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23896\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__23899\,
            I => \buf_readRTD_11\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23896\,
            I => \buf_readRTD_11\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__23885\,
            I => n22214
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23876\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23872\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__23875\,
            I => \N__23869\
        );

    \I__3134\ : Span4Mux_h
    port map (
            O => \N__23872\,
            I => \N__23866\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23863\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__23866\,
            I => buf_adcdata_vdc_19
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23863\,
            I => buf_adcdata_vdc_19
        );

    \I__3130\ : InMux
    port map (
            O => \N__23858\,
            I => \N__23855\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__23855\,
            I => \N__23851\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23848\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__23851\,
            I => \N__23845\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23848\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__23845\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23837\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__23837\,
            I => \N__23833\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23830\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__23833\,
            I => \N__23827\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23830\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__23827\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23812\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23809\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__23812\,
            I => \N__23806\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__23809\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__23806\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23794\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23791\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__23794\,
            I => \N__23788\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23791\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__23788\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23777\
        );

    \I__3103\ : Odrv12
    port map (
            O => \N__23777\,
            I => \ADC_VDC.n21\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__23774\,
            I => \n12875_cascade_\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23763\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23758\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23758\
        );

    \I__3097\ : Span12Mux_s9_v
    port map (
            O => \N__23763\,
            I => \N__23755\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23758\,
            I => buf_adcdata_iac_6
        );

    \I__3095\ : Odrv12
    port map (
            O => \N__23755\,
            I => buf_adcdata_iac_6
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__23750\,
            I => \n19_adj_1628_cascade_\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23741\
        );

    \I__3091\ : Span12Mux_h
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__3090\ : Odrv12
    port map (
            O => \N__23738\,
            I => buf_data_iac_6
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__23735\,
            I => \n22_adj_1629_cascade_\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23732\,
            I => \N__23728\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23720\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23728\,
            I => \N__23720\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23720\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__23720\,
            I => cmd_rdadctmp_14_adj_1436
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__23717\,
            I => \N__23713\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__23716\,
            I => \N__23710\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23706\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23701\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23701\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23706\,
            I => cmd_rdadctmp_15_adj_1435
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23701\,
            I => cmd_rdadctmp_15_adj_1435
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__23696\,
            I => \N__23692\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23687\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23687\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23683\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23680\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__23683\,
            I => cmd_rdadctmp_14
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__23680\,
            I => cmd_rdadctmp_14
        );

    \I__3069\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23672\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__23672\,
            I => \N__23668\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__23671\,
            I => \N__23665\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__23668\,
            I => \N__23662\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23659\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__23662\,
            I => buf_adcdata_vdc_7
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__23659\,
            I => buf_adcdata_vdc_7
        );

    \I__3062\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23647\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23643\
        );

    \I__3059\ : Span4Mux_h
    port map (
            O => \N__23647\,
            I => \N__23640\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23637\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__23643\,
            I => buf_adcdata_vac_7
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__23640\,
            I => buf_adcdata_vac_7
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23637\,
            I => buf_adcdata_vac_7
        );

    \I__3054\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__3052\ : Span12Mux_s8_v
    port map (
            O => \N__23624\,
            I => \N__23619\
        );

    \I__3051\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23614\
        );

    \I__3050\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23614\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__23619\,
            I => buf_adcdata_iac_7
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__23614\,
            I => buf_adcdata_iac_7
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__23609\,
            I => \n19_adj_1625_cascade_\
        );

    \I__3046\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__3044\ : Span12Mux_h
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__3043\ : Odrv12
    port map (
            O => \N__23597\,
            I => buf_data_iac_7
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__23594\,
            I => \n22_adj_1626_cascade_\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23587\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__23590\,
            I => \N__23584\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23587\,
            I => \N__23580\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23577\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23574\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__23580\,
            I => \N__23571\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__23577\,
            I => buf_adcdata_vac_6
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__23574\,
            I => buf_adcdata_vac_6
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__23571\,
            I => buf_adcdata_vac_6
        );

    \I__3032\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__23558\,
            I => \N__23554\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23551\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__23554\,
            I => buf_adcdata_vdc_6
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__23551\,
            I => buf_adcdata_vdc_6
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23540\,
            I => \CLK_DDS.tmp_buf_14\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23530\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23527\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23524\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__23527\,
            I => \N__23519\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__23524\,
            I => \N__23519\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__23516\,
            I => tmp_buf_15_adj_1455
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__23513\,
            I => \N__23500\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__23512\,
            I => \N__23491\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23485\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23480\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23465\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23465\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23465\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23465\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23465\
        );

    \I__3006\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23465\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23465\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23460\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23460\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23451\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23451\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23451\
        );

    \I__2999\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23451\
        );

    \I__2998\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23444\
        );

    \I__2997\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23444\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23444\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23441\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23437\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23485\,
            I => \N__23434\
        );

    \I__2992\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23431\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23428\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23425\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23422\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23412\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23412\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23412\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23412\
        );

    \I__2984\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23409\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23406\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__23434\,
            I => \N__23403\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23394\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23428\,
            I => \N__23394\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__23425\,
            I => \N__23394\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__23422\,
            I => \N__23394\
        );

    \I__2977\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23389\
        );

    \I__2976\ : Span4Mux_v
    port map (
            O => \N__23412\,
            I => \N__23386\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23377\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__23406\,
            I => \N__23377\
        );

    \I__2973\ : Span4Mux_v
    port map (
            O => \N__23403\,
            I => \N__23377\
        );

    \I__2972\ : Span4Mux_v
    port map (
            O => \N__23394\,
            I => \N__23377\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23372\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23372\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__23389\,
            I => \N__23367\
        );

    \I__2968\ : Span4Mux_h
    port map (
            O => \N__23386\,
            I => \N__23367\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__23377\,
            I => dds_state_2_adj_1452
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__23372\,
            I => dds_state_2_adj_1452
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__23367\,
            I => dds_state_2_adj_1452
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__2963\ : SRMux
    port map (
            O => \N__23359\,
            I => \N__23349\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23346\
        );

    \I__2961\ : CEMux
    port map (
            O => \N__23357\,
            I => \N__23343\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23328\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__23353\,
            I => \N__23320\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23313\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23310\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23305\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23343\,
            I => \N__23305\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23302\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23287\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23287\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23287\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23287\
        );

    \I__2949\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23287\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23287\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23287\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23334\,
            I => \N__23278\
        );

    \I__2945\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23278\
        );

    \I__2944\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23278\
        );

    \I__2943\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23278\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23328\,
            I => \N__23275\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23264\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23264\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23264\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23264\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23264\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23261\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23258\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23255\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23317\,
            I => \N__23252\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23316\,
            I => \N__23249\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23246\
        );

    \I__2930\ : Span4Mux_h
    port map (
            O => \N__23310\,
            I => \N__23243\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__23305\,
            I => \N__23240\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__23302\,
            I => \N__23229\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23229\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__23278\,
            I => \N__23229\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__23275\,
            I => \N__23229\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23264\,
            I => \N__23229\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23217\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23217\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23255\,
            I => \N__23217\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__23252\,
            I => \N__23217\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__23249\,
            I => \N__23217\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__23246\,
            I => \N__23214\
        );

    \I__2917\ : Span4Mux_h
    port map (
            O => \N__23243\,
            I => \N__23207\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23207\
        );

    \I__2915\ : Span4Mux_v
    port map (
            O => \N__23229\,
            I => \N__23207\
        );

    \I__2914\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23204\
        );

    \I__2913\ : Odrv12
    port map (
            O => \N__23217\,
            I => dds_state_1_adj_1453
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__23214\,
            I => dds_state_1_adj_1453
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__23207\,
            I => dds_state_1_adj_1453
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23204\,
            I => dds_state_1_adj_1453
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23189\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__23189\,
            I => \CLK_DDS.tmp_buf_8\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__2905\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23180\,
            I => \CLK_DDS.tmp_buf_9\
        );

    \I__2903\ : CEMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__23171\,
            I => \N__23166\
        );

    \I__2900\ : CEMux
    port map (
            O => \N__23170\,
            I => \N__23163\
        );

    \I__2899\ : CEMux
    port map (
            O => \N__23169\,
            I => \N__23160\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__23166\,
            I => \N__23155\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23155\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23152\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23149\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__23152\,
            I => \N__23146\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__23149\,
            I => \N__23139\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__23146\,
            I => \N__23139\
        );

    \I__2891\ : CEMux
    port map (
            O => \N__23145\,
            I => \N__23136\
        );

    \I__2890\ : CEMux
    port map (
            O => \N__23144\,
            I => \N__23133\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__23139\,
            I => \CLK_DDS.n12800\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__23136\,
            I => \CLK_DDS.n12800\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__23133\,
            I => \CLK_DDS.n12800\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__23126\,
            I => \N__23122\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__23125\,
            I => \N__23118\
        );

    \I__2884\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23115\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__23121\,
            I => \N__23111\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23108\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__23115\,
            I => \N__23105\
        );

    \I__2880\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23100\
        );

    \I__2879\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23100\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__23108\,
            I => trig_dds1
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__23105\,
            I => trig_dds1
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__23100\,
            I => trig_dds1
        );

    \I__2875\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23090\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__2873\ : Span4Mux_v
    port map (
            O => \N__23087\,
            I => \N__23084\
        );

    \I__2872\ : Sp12to4
    port map (
            O => \N__23084\,
            I => \N__23081\
        );

    \I__2871\ : Span12Mux_h
    port map (
            O => \N__23081\,
            I => \N__23078\
        );

    \I__2870\ : Odrv12
    port map (
            O => \N__23078\,
            I => \ICE_GPMO_1\
        );

    \I__2869\ : IoInMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__2867\ : IoSpan4Mux
    port map (
            O => \N__23069\,
            I => \N__23065\
        );

    \I__2866\ : IoInMux
    port map (
            O => \N__23068\,
            I => \N__23062\
        );

    \I__2865\ : IoSpan4Mux
    port map (
            O => \N__23065\,
            I => \N__23059\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__23056\
        );

    \I__2863\ : Span4Mux_s2_v
    port map (
            O => \N__23059\,
            I => \N__23053\
        );

    \I__2862\ : IoSpan4Mux
    port map (
            O => \N__23056\,
            I => \N__23050\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__23053\,
            I => \N__23047\
        );

    \I__2860\ : Sp12to4
    port map (
            O => \N__23050\,
            I => \N__23044\
        );

    \I__2859\ : Sp12to4
    port map (
            O => \N__23047\,
            I => \N__23039\
        );

    \I__2858\ : Span12Mux_h
    port map (
            O => \N__23044\,
            I => \N__23039\
        );

    \I__2857\ : Span12Mux_v
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__23036\,
            I => \IAC_CLK\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__2854\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__23027\,
            I => n22100
        );

    \I__2852\ : IoInMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__23018\
        );

    \I__2850\ : IoSpan4Mux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__2849\ : Span4Mux_s0_v
    port map (
            O => \N__23015\,
            I => \N__23012\
        );

    \I__2848\ : Sp12to4
    port map (
            O => \N__23012\,
            I => \N__23008\
        );

    \I__2847\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23004\
        );

    \I__2846\ : Span12Mux_v
    port map (
            O => \N__23008\,
            I => \N__23001\
        );

    \I__2845\ : InMux
    port map (
            O => \N__23007\,
            I => \N__22998\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__22995\
        );

    \I__2843\ : Odrv12
    port map (
            O => \N__23001\,
            I => \SELIRNG0\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__22998\,
            I => \SELIRNG0\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__22995\,
            I => \SELIRNG0\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22982\,
            I => \CLK_DDS.tmp_buf_10\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__22979\,
            I => \N__22976\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22973\,
            I => \CLK_DDS.tmp_buf_11\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22964\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22964\,
            I => \CLK_DDS.tmp_buf_12\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22958\,
            I => \CLK_DDS.tmp_buf_13\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__22955\,
            I => \N__22951\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22947\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22944\
        );

    \I__2826\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22941\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22938\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__22944\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22941\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22938\,
            I => cmd_rdadctmp_25_adj_1425
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__22931\,
            I => \N__22927\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__22930\,
            I => \N__22924\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22921\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22918\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22921\,
            I => cmd_rdadctmp_31_adj_1419
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22918\,
            I => cmd_rdadctmp_31_adj_1419
        );

    \I__2815\ : IoInMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__2813\ : Span12Mux_s11_h
    port map (
            O => \N__22907\,
            I => \N__22902\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22897\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22897\
        );

    \I__2810\ : Odrv12
    port map (
            O => \N__22902\,
            I => \VAC_OSR1\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22897\,
            I => \VAC_OSR1\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22886\
        );

    \I__2806\ : Span4Mux_v
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__2805\ : Sp12to4
    port map (
            O => \N__22883\,
            I => \N__22878\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__22882\,
            I => \N__22875\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22872\
        );

    \I__2802\ : Span12Mux_h
    port map (
            O => \N__22878\,
            I => \N__22869\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22866\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__22872\,
            I => buf_adcdata_iac_21
        );

    \I__2799\ : Odrv12
    port map (
            O => \N__22869\,
            I => buf_adcdata_iac_21
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__22866\,
            I => buf_adcdata_iac_21
        );

    \I__2797\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__2795\ : Span12Mux_h
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__2794\ : Span12Mux_v
    port map (
            O => \N__22850\,
            I => \N__22845\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22840\
        );

    \I__2792\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22840\
        );

    \I__2791\ : Odrv12
    port map (
            O => \N__22845\,
            I => buf_adcdata_iac_23
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__22840\,
            I => buf_adcdata_iac_23
        );

    \I__2789\ : IoInMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22832\,
            I => \N__22829\
        );

    \I__2787\ : IoSpan4Mux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__2786\ : Span4Mux_s0_h
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__2785\ : Sp12to4
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__2784\ : Span12Mux_s11_h
    port map (
            O => \N__22820\,
            I => \N__22815\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22810\
        );

    \I__2782\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22810\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__22815\,
            I => \VAC_FLT1\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22810\,
            I => \VAC_FLT1\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__2777\ : Span4Mux_v
    port map (
            O => \N__22799\,
            I => \N__22796\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__22796\,
            I => n17_adj_1525
        );

    \I__2775\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22790\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__22790\,
            I => \N__22787\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__2772\ : Sp12to4
    port map (
            O => \N__22784\,
            I => \N__22779\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22776\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22773\
        );

    \I__2769\ : Span12Mux_h
    port map (
            O => \N__22779\,
            I => \N__22770\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22767\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22773\,
            I => buf_adcdata_iac_16
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__22770\,
            I => buf_adcdata_iac_16
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22767\,
            I => buf_adcdata_iac_16
        );

    \I__2764\ : IoInMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__2762\ : Span4Mux_s2_v
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__2759\ : Sp12to4
    port map (
            O => \N__22745\,
            I => \N__22740\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22735\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22735\
        );

    \I__2756\ : Odrv12
    port map (
            O => \N__22740\,
            I => \IAC_OSR0\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22735\,
            I => \IAC_OSR0\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__22730\,
            I => \RTD.n21276_cascade_\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22724\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22724\,
            I => \RTD.n21275\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22717\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22714\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22717\,
            I => \RTD.adc_state_3_N_1368_1\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__22714\,
            I => \RTD.adc_state_3_N_1368_1\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \RTD.adc_state_3_N_1368_1_cascade_\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22703\,
            I => \RTD.n7\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__2743\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__22688\,
            I => \RTD.n20762\
        );

    \I__2739\ : CEMux
    port map (
            O => \N__22685\,
            I => \N__22680\
        );

    \I__2738\ : CEMux
    port map (
            O => \N__22684\,
            I => \N__22677\
        );

    \I__2737\ : CEMux
    port map (
            O => \N__22683\,
            I => \N__22674\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22671\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__22677\,
            I => \N__22668\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22665\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__22671\,
            I => \RTD.n11742\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__22668\,
            I => \RTD.n11742\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__22665\,
            I => \RTD.n11742\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__22658\,
            I => \n16_adj_1512_cascade_\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__22655\,
            I => \RTD.n21323_cascade_\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__22649\,
            I => \RTD.n26\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__22646\,
            I => \RTD.n21325_cascade_\
        );

    \I__2725\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22640\,
            I => \RTD.n4\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22634\,
            I => \N__22629\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22624\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22624\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__22629\,
            I => \RTD.n1\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__22624\,
            I => \RTD.n1\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__22619\,
            I => \RTD.n1_cascade_\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22609\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__22612\,
            I => \RTD.n20587\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22609\,
            I => \RTD.n20587\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__22598\,
            I => n8_adj_1608
        );

    \I__2709\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__2707\ : Span4Mux_v
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__2706\ : Odrv4
    port map (
            O => \N__22586\,
            I => n21227
        );

    \I__2705\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22577\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22570\
        );

    \I__2703\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22567\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22564\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22561\
        );

    \I__2700\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22556\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22556\
        );

    \I__2698\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22553\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22550\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__22570\,
            I => \N__22547\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22567\,
            I => \N__22544\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22564\,
            I => \N__22540\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__22561\,
            I => \N__22533\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22533\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22533\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22550\,
            I => \N__22529\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__22547\,
            I => \N__22524\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__22544\,
            I => \N__22524\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22521\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__22540\,
            I => \N__22516\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__22533\,
            I => \N__22516\
        );

    \I__2684\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22513\
        );

    \I__2683\ : Span4Mux_h
    port map (
            O => \N__22529\,
            I => \N__22508\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__22524\,
            I => \N__22508\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22505\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__22516\,
            I => \N__22502\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22513\,
            I => dds_state_0_adj_1454
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__22508\,
            I => dds_state_0_adj_1454
        );

    \I__2677\ : Odrv12
    port map (
            O => \N__22505\,
            I => dds_state_0_adj_1454
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__22502\,
            I => dds_state_0_adj_1454
        );

    \I__2675\ : CEMux
    port map (
            O => \N__22493\,
            I => \N__22489\
        );

    \I__2674\ : CEMux
    port map (
            O => \N__22492\,
            I => \N__22486\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__22489\,
            I => \N__22483\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22480\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__22483\,
            I => \N__22477\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__22480\,
            I => \N__22474\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__22477\,
            I => \CLK_DDS.n9\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__22474\,
            I => \CLK_DDS.n9\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__22469\,
            I => \N__22465\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__22468\,
            I => \N__22462\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22458\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22455\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__22461\,
            I => \N__22451\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22448\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__22455\,
            I => \N__22445\
        );

    \I__2660\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22440\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22440\
        );

    \I__2658\ : Span4Mux_h
    port map (
            O => \N__22448\,
            I => \N__22437\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__22445\,
            I => \RTD.mode\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__22440\,
            I => \RTD.mode\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__22437\,
            I => \RTD.mode\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22422\
        );

    \I__2652\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22417\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22417\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__22422\,
            I => \N__22412\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22412\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__2646\ : Sp12to4
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2645\ : Span12Mux_v
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__22400\,
            I => \RTD_DRDY\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__2641\ : Span4Mux_h
    port map (
            O => \N__22391\,
            I => \N__22384\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22379\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22379\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22376\
        );

    \I__2637\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22373\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__22384\,
            I => \RTD.adress_7_N_1340_7\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__22379\,
            I => \RTD.adress_7_N_1340_7\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22376\,
            I => \RTD.adress_7_N_1340_7\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22373\,
            I => \RTD.adress_7_N_1340_7\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__22361\,
            I => \RTD.n16669\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \RTD.n16669_cascade_\
        );

    \I__2629\ : IoInMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2627\ : IoSpan4Mux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2626\ : Span4Mux_s0_h
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2625\ : Sp12to4
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2624\ : Span12Mux_s11_h
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__2623\ : Odrv12
    port map (
            O => \N__22337\,
            I => \RTD_CS\
        );

    \I__2622\ : CEMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__22319\,
            I => \RTD.n11703\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22312\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22309\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22312\,
            I => \RTD.cfg_buf_1\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22309\,
            I => \RTD.cfg_buf_1\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__22301\,
            I => \RTD.n12_adj_1397\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22291\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__2607\ : Span4Mux_h
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22282\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__22285\,
            I => buf_adcdata_vdc_23
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__22282\,
            I => buf_adcdata_vdc_23
        );

    \I__2603\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__2599\ : Sp12to4
    port map (
            O => \N__22265\,
            I => \N__22260\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22257\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22254\
        );

    \I__2596\ : Span12Mux_h
    port map (
            O => \N__22260\,
            I => \N__22249\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22249\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__22254\,
            I => buf_adcdata_vac_23
        );

    \I__2593\ : Odrv12
    port map (
            O => \N__22249\,
            I => buf_adcdata_vac_23
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__22244\,
            I => \n19_adj_1526_cascade_\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__22241\,
            I => \n22076_cascade_\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__22232\,
            I => \N__22228\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22225\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__22228\,
            I => \buf_readRTD_15\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__22225\,
            I => \buf_readRTD_15\
        );

    \I__2584\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__22217\,
            I => n20
        );

    \I__2582\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__22208\,
            I => \RTD.n22370\
        );

    \I__2579\ : IoInMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2577\ : IoSpan4Mux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__2576\ : Span4Mux_s3_h
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2575\ : Span4Mux_h
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2573\ : Sp12to4
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__22184\,
            I => \RTD_SCLK\
        );

    \I__2571\ : CEMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__22172\,
            I => \RTD.n8\
        );

    \I__2567\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22147\
        );

    \I__2566\ : InMux
    port map (
            O => \N__22168\,
            I => \N__22147\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22147\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22140\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22140\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22140\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22133\
        );

    \I__2560\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22133\
        );

    \I__2559\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22133\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22118\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22118\
        );

    \I__2556\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22118\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22118\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22118\
        );

    \I__2553\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22118\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22118\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22115\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22112\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__22133\,
            I => \N__22109\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22106\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__22115\,
            I => \N__22103\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__22112\,
            I => \N__22098\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__22109\,
            I => \N__22098\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__22106\,
            I => \N__22095\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__22103\,
            I => n13309
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__22098\,
            I => n13309
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__22095\,
            I => n13309
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__22088\,
            I => \N__22083\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22076\
        );

    \I__2538\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22076\
        );

    \I__2537\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22076\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__22076\,
            I => cmd_rdadctmp_30
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \N__22069\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__22072\,
            I => \N__22066\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22061\
        );

    \I__2532\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22061\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__22061\,
            I => cmd_rdadctmp_31
        );

    \I__2530\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__22051\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22048\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__22051\,
            I => buf_adcdata_vdc_5
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__22048\,
            I => buf_adcdata_vdc_5
        );

    \I__2525\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__22040\,
            I => \N__22036\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22033\
        );

    \I__2522\ : Odrv12
    port map (
            O => \N__22036\,
            I => buf_adcdata_vdc_4
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__22033\,
            I => buf_adcdata_vdc_4
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__2519\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__22022\,
            I => \N__22018\
        );

    \I__2517\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22015\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__22018\,
            I => buf_adcdata_vdc_20
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__22015\,
            I => buf_adcdata_vdc_20
        );

    \I__2514\ : CEMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__22001\,
            I => \ADC_VDC.n47\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21986\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21986\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21986\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21986\,
            I => cmd_rdadctmp_15
        );

    \I__2505\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21980\,
            I => n19_adj_1631
        );

    \I__2503\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21970\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21966\
        );

    \I__2500\ : Span12Mux_s10_v
    port map (
            O => \N__21970\,
            I => \N__21963\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21960\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21966\,
            I => buf_adcdata_vac_5
        );

    \I__2497\ : Odrv12
    port map (
            O => \N__21963\,
            I => buf_adcdata_vac_5
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__21960\,
            I => buf_adcdata_vac_5
        );

    \I__2495\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2492\ : Sp12to4
    port map (
            O => \N__21944\,
            I => \N__21939\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21936\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21933\
        );

    \I__2489\ : Span12Mux_h
    port map (
            O => \N__21939\,
            I => \N__21928\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21928\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21933\,
            I => buf_adcdata_vac_20
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__21928\,
            I => buf_adcdata_vac_20
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \N__21919\
        );

    \I__2484\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21916\,
            I => \N__21910\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21913\,
            I => \N__21906\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__21910\,
            I => \N__21903\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21900\
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__21906\,
            I => cmd_rdadctmp_29
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__21903\,
            I => cmd_rdadctmp_29
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__21900\,
            I => cmd_rdadctmp_29
        );

    \I__2475\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__21887\,
            I => \N__21882\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21877\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21877\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__21882\,
            I => buf_adcdata_vac_4
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21877\,
            I => buf_adcdata_vac_4
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21872\,
            I => \n19_adj_1636_cascade_\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__21863\,
            I => \N__21858\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21853\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21853\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__21858\,
            I => buf_adcdata_iac_4
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21853\,
            I => buf_adcdata_iac_4
        );

    \I__2460\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__21839\,
            I => buf_data_iac_4
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__21836\,
            I => \n22_adj_1637_cascade_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21827\
        );

    \I__2453\ : Span12Mux_v
    port map (
            O => \N__21827\,
            I => \N__21823\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21820\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__21823\,
            I => cmd_rdadctmp_4
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21820\,
            I => cmd_rdadctmp_4
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__21815\,
            I => \N__21811\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21806\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21806\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21806\,
            I => cmd_rdadctmp_5
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21797\,
            I => \CLK_DDS.tmp_buf_2\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21788\,
            I => \CLK_DDS.tmp_buf_3\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21779\,
            I => \CLK_DDS.tmp_buf_4\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21773\,
            I => \CLK_DDS.tmp_buf_5\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2433\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21764\,
            I => \CLK_DDS.tmp_buf_6\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21758\,
            I => \CLK_DDS.tmp_buf_7\
        );

    \I__2429\ : CEMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__21743\,
            I => \CLK_DDS.n9_adj_1395\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21730\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21730\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21727\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21730\,
            I => cmd_rdadctmp_30_adj_1420
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__21727\,
            I => cmd_rdadctmp_30_adj_1420
        );

    \I__2418\ : IoInMux
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__2416\ : Span12Mux_s9_v
    port map (
            O => \N__21716\,
            I => \N__21712\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__2414\ : Odrv12
    port map (
            O => \N__21712\,
            I => \DDS_MOSI1\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21709\,
            I => \DDS_MOSI1\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21696\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21691\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21691\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__21696\,
            I => cmd_rdadctmp_23_adj_1427
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__21691\,
            I => cmd_rdadctmp_23_adj_1427
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__21686\,
            I => \N__21682\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__21685\,
            I => \N__21678\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21671\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21671\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21671\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21671\,
            I => cmd_rdadctmp_24_adj_1426
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__21668\,
            I => \N__21663\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__21667\,
            I => \N__21660\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21655\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21655\
        );

    \I__2396\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21652\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__21655\,
            I => cmd_rdadctmp_26_adj_1424
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__21652\,
            I => cmd_rdadctmp_26_adj_1424
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__2392\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__21632\,
            I => \CLK_DDS.tmp_buf_1\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__21629\,
            I => \N__21625\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21618\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21613\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21613\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21618\,
            I => read_buf_7
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__21613\,
            I => read_buf_7
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__21608\,
            I => \N__21603\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__21607\,
            I => \N__21600\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21595\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21595\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21592\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21595\,
            I => read_buf_2
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21592\,
            I => read_buf_2
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__21587\,
            I => \N__21582\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__21586\,
            I => \N__21579\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__21585\,
            I => \N__21576\
        );

    \I__2370\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21573\
        );

    \I__2369\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21568\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21568\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__21573\,
            I => read_buf_3
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__21568\,
            I => read_buf_3
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__21563\,
            I => \N__21556\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__21561\,
            I => \N__21550\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__21560\,
            I => \N__21547\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__21559\,
            I => \N__21542\
        );

    \I__2360\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21529\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21529\
        );

    \I__2358\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21529\
        );

    \I__2357\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21529\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21529\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21529\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21526\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21513\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21513\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21510\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21505\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21505\
        );

    \I__2348\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21498\
        );

    \I__2347\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21498\
        );

    \I__2346\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21498\
        );

    \I__2345\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21493\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21493\
        );

    \I__2343\ : Span4Mux_h
    port map (
            O => \N__21513\,
            I => \N__21490\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__21510\,
            I => n1_adj_1601
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21505\,
            I => n1_adj_1601
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21498\,
            I => n1_adj_1601
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__21493\,
            I => n1_adj_1601
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__21490\,
            I => n1_adj_1601
        );

    \I__2337\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21470\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21470\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21470\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21470\,
            I => read_buf_4
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__21467\,
            I => \n1_adj_1601_cascade_\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21459\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21454\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21454\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__21459\,
            I => read_buf_5
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__21454\,
            I => read_buf_5
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \N__21445\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__21448\,
            I => \N__21441\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21438\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21433\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21433\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__21438\,
            I => cmd_rdadctmp_29_adj_1421
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21433\,
            I => cmd_rdadctmp_29_adj_1421
        );

    \I__2320\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21425\,
            I => \RTD.cfg_tmp_2\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21419\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21419\,
            I => \RTD.cfg_tmp_3\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21413\,
            I => \RTD.cfg_tmp_4\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21407\,
            I => \RTD.cfg_tmp_5\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21401\,
            I => \RTD.cfg_tmp_6\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21391\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21388\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__21391\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21388\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2305\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__21380\,
            I => \RTD.cfg_tmp_0\
        );

    \I__2303\ : CEMux
    port map (
            O => \N__21377\,
            I => \N__21373\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21370\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__21373\,
            I => \RTD.n13228\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21370\,
            I => \RTD.n13228\
        );

    \I__2299\ : SRMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__21356\,
            I => \RTD.n15015\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__21353\,
            I => \RTD.n7333_cascade_\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \RTD.n13_cascade_\
        );

    \I__2293\ : CEMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__21341\,
            I => \RTD.n11734\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21330\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21327\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21324\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__21330\,
            I => \RTD.n7333\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__21327\,
            I => \RTD.n7333\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21324\,
            I => \RTD.n7333\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21314\,
            I => \RTD.cfg_tmp_1\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21308\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21295\
        );

    \I__2276\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__21295\,
            I => read_buf_15
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21292\,
            I => read_buf_15
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__21287\,
            I => \n11730_cascade_\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21280\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21277\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21280\,
            I => adress_6
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__21277\,
            I => adress_6
        );

    \I__2268\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21268\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21265\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21268\,
            I => \RTD.cfg_buf_6\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21265\,
            I => \RTD.cfg_buf_6\
        );

    \I__2264\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21256\
        );

    \I__2263\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21253\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__21256\,
            I => \RTD.cfg_buf_0\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__21253\,
            I => \RTD.cfg_buf_0\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__21248\,
            I => \RTD.n9_cascade_\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__21245\,
            I => \RTD.adress_7_N_1340_7_cascade_\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21235\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21232\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21235\,
            I => \RTD.adress_7\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21232\,
            I => \RTD.adress_7\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__2252\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__21218\,
            I => adress_0
        );

    \I__2249\ : CEMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21203\
        );

    \I__2247\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21192\
        );

    \I__2246\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21192\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21192\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21192\
        );

    \I__2243\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21192\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21189\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__21203\,
            I => n13181
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__21192\,
            I => n13181
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__21189\,
            I => n13181
        );

    \I__2238\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21178\
        );

    \I__2237\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21175\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__21178\,
            I => \RTD.cfg_buf_5\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__21175\,
            I => \RTD.cfg_buf_5\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__2233\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21163\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21160\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__21163\,
            I => \RTD.cfg_buf_3\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21160\,
            I => \RTD.cfg_buf_3\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__21152\,
            I => \RTD.n11\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \ADC_VDC.n13038_cascade_\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__21140\,
            I => \ADC_VDC.n20659\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__21137\,
            I => \ADC_VDC.n17432_cascade_\
        );

    \I__2222\ : SRMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__21125\,
            I => \ADC_VDC.n18466\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__2217\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21112\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__21115\,
            I => \N__21108\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__21112\,
            I => \N__21105\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21100\
        );

    \I__2212\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21100\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__21105\,
            I => read_buf_11
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__21100\,
            I => read_buf_11
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \ADC_VDC.n11692_cascade_\
        );

    \I__2208\ : IoInMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__21089\,
            I => \N__21085\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21082\
        );

    \I__2205\ : Span12Mux_s5_h
    port map (
            O => \N__21085\,
            I => \N__21079\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21076\
        );

    \I__2203\ : Odrv12
    port map (
            O => \N__21079\,
            I => \VDC_SCLK\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__21076\,
            I => \VDC_SCLK\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__21071\,
            I => \N__21064\
        );

    \I__2200\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21061\
        );

    \I__2199\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21058\
        );

    \I__2198\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21053\
        );

    \I__2197\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21053\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21050\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__21061\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__21058\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__21053\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__21050\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__2191\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21037\
        );

    \I__2190\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21034\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__21037\,
            I => \ADC_VDC.n20534\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__21034\,
            I => \ADC_VDC.n20534\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__21029\,
            I => \N__21024\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__21028\,
            I => \N__21021\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__21027\,
            I => \N__21017\
        );

    \I__2184\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21011\
        );

    \I__2183\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21011\
        );

    \I__2182\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21008\
        );

    \I__2181\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21005\
        );

    \I__2180\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21002\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__20999\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__21008\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__21005\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__21002\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__20999\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__20981\,
            I => \ADC_VDC.n6_adj_1410\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__20978\,
            I => \ADC_VDC.n11281_cascade_\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20968\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20965\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20960\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20960\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20957\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20968\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20965\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20960\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__20957\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20942\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20942\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20942\,
            I => \ADC_VDC.n15\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__20939\,
            I => \ADC_VDC.n15_cascade_\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__20936\,
            I => \ADC_VDC.n20746_cascade_\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20930\,
            I => \ADC_VDC.n72\
        );

    \I__2153\ : CEMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__20921\,
            I => \ADC_VDC.n12823\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__20918\,
            I => \ADC_VDC.n19_adj_1413_cascade_\
        );

    \I__2149\ : CEMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20912\,
            I => \ADC_VDC.n17\
        );

    \I__2147\ : SRMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__20900\,
            I => \ADC_VDC.n4\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__20897\,
            I => \ADC_VDC.n10132_cascade_\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20888\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20888\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20888\,
            I => \ADC_VDC.n7_adj_1411\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20879\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20879\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__20879\,
            I => \ADC_VDC.n20750\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20873\,
            I => \ADC_VDC.n12\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__20870\,
            I => \ADC_VDC.n20750_cascade_\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20863\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20863\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20860\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20855\,
            I => \ADC_IAC.n19418\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20848\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20845\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__20848\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20845\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20840\,
            I => \ADC_IAC.n19419\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20833\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20830\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__20833\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20830\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20825\,
            I => \ADC_IAC.n19420\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20822\,
            I => \ADC_IAC.n19421\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20815\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20812\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__20815\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__20812\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__2113\ : CEMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__2110\ : Span4Mux_h
    port map (
            O => \N__20798\,
            I => \N__20794\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20791\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__20794\,
            I => \ADC_IAC.n12586\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20791\,
            I => \ADC_IAC.n12586\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__20786\,
            I => \N__20783\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2104\ : Span4Mux_h
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__20777\,
            I => \ADC_IAC.n14860\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \N__20770\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20764\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20767\,
            I => cmd_rdadctmp_1_adj_1449
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__20764\,
            I => cmd_rdadctmp_1_adj_1449
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20752\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \N__20749\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20752\,
            I => \N__20746\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__20746\,
            I => cmd_rdadctmp_2_adj_1448
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20743\,
            I => cmd_rdadctmp_2_adj_1448
        );

    \I__2090\ : IoInMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__2088\ : Span4Mux_s2_v
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__20723\,
            I => \DDS_MCLK1\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__20711\,
            I => \N__20707\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__20710\,
            I => \N__20703\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__20707\,
            I => \N__20700\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20697\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20694\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__20700\,
            I => cmd_rdadctmp_28_adj_1422
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20697\,
            I => cmd_rdadctmp_28_adj_1422
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__20694\,
            I => cmd_rdadctmp_28_adj_1422
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20678\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20678\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__20678\,
            I => cmd_rdadctmp_3_adj_1447
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20666\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20663\
        );

    \I__2066\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20658\
        );

    \I__2065\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20658\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20650\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20663\,
            I => \N__20650\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20650\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__20657\,
            I => \N__20647\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__20650\,
            I => \N__20644\
        );

    \I__2059\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20641\
        );

    \I__2058\ : Sp12to4
    port map (
            O => \N__20644\,
            I => \N__20636\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__20641\,
            I => \N__20636\
        );

    \I__2056\ : Span12Mux_h
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__2055\ : Odrv12
    port map (
            O => \N__20633\,
            I => \IAC_DRDY\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20627\,
            I => n20612
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__20624\,
            I => \n14_adj_1604_cascade_\
        );

    \I__2051\ : IoInMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20618\,
            I => \N__20615\
        );

    \I__2049\ : IoSpan4Mux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2048\ : Sp12to4
    port map (
            O => \N__20612\,
            I => \N__20608\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__20611\,
            I => \N__20605\
        );

    \I__2046\ : Span12Mux_v
    port map (
            O => \N__20608\,
            I => \N__20602\
        );

    \I__2045\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20599\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__20602\,
            I => \IAC_CS\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__20599\,
            I => \IAC_CS\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20590\
        );

    \I__2041\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__20590\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__20587\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20582\,
            I => \bfn_6_15_0_\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__20579\,
            I => \N__20575\
        );

    \I__2036\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20569\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20572\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__20569\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__2032\ : InMux
    port map (
            O => \N__20564\,
            I => \ADC_IAC.n19415\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20557\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20554\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20557\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20554\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20549\,
            I => \ADC_IAC.n19416\
        );

    \I__2026\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20542\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20539\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20542\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__20539\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__2022\ : InMux
    port map (
            O => \N__20534\,
            I => \ADC_IAC.n19417\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20520\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20515\
        );

    \I__2017\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20515\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__20520\,
            I => read_buf_13
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20515\,
            I => read_buf_13
        );

    \I__2014\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20507\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__20507\,
            I => \N__20502\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20497\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20497\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__20502\,
            I => read_buf_8
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__20497\,
            I => read_buf_8
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__20492\,
            I => \N__20487\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__20491\,
            I => \N__20483\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20471\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20471\
        );

    \I__2004\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20471\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20471\
        );

    \I__2002\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20471\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__20471\,
            I => \N__20467\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__1999\ : Odrv12
    port map (
            O => \N__20467\,
            I => n20754
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__20464\,
            I => n20754
        );

    \I__1997\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20455\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__20455\,
            I => cmd_rdadctmp_5_adj_1445
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20452\,
            I => cmd_rdadctmp_5_adj_1445
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20438\
        );

    \I__1991\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20438\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__20438\,
            I => cmd_rdadctmp_4_adj_1446
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__20435\,
            I => \RTD.n19_cascade_\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__20432\,
            I => \N__20427\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20424\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20419\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20419\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20424\,
            I => read_buf_9
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__20419\,
            I => read_buf_9
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__1981\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__20408\,
            I => \N__20404\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__20404\,
            I => adress_1
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__20401\,
            I => adress_1
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20391\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \N__20388\
        );

    \I__1974\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20381\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20381\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20381\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20381\,
            I => read_buf_1
        );

    \I__1970\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20372\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20372\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__20372\,
            I => adress_2
        );

    \I__1967\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20363\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20363\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__20363\,
            I => adress_4
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20351\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20351\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20351\,
            I => adress_5
        );

    \I__1960\ : IoInMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__1958\ : Span4Mux_s1_h
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__1956\ : Span4Mux_v
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__20327\,
            I => \RTD_SDI\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \RTD.n21309_cascade_\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__20318\,
            I => \RTD.n12\
        );

    \I__1949\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20311\
        );

    \I__1948\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20305\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__20311\,
            I => \N__20302\
        );

    \I__1946\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20299\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20294\
        );

    \I__1944\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20294\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__20305\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__20302\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__20299\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__20294\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__20282\,
            I => \ADC_VDC.n6\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__20279\,
            I => \ADC_VDC.n10552_cascade_\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__20273\,
            I => \ADC_VDC.n21974\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20262\
        );

    \I__1933\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20262\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__20268\,
            I => \N__20259\
        );

    \I__1931\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20255\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__20262\,
            I => \N__20252\
        );

    \I__1929\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20249\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20246\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__20255\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__20252\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20249\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20246\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__20231\,
            I => \ADC_VDC.n20562\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20228\,
            I => \ADC_VDC.n21224_cascade_\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__20219\,
            I => \ADC_VDC.n20748\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__20216\,
            I => \ADC_VDC.n31_cascade_\
        );

    \I__1915\ : CEMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__20204\,
            I => \ADC_VDC.n20555\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20193\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20188\
        );

    \I__1908\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20188\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__20193\,
            I => read_buf_12
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20188\,
            I => read_buf_12
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__1904\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20174\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20174\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__20174\,
            I => adress_3
        );

    \I__1901\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20166\
        );

    \I__1900\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20163\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20160\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20166\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__20163\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__20160\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \ADC_VDC.n20534_cascade_\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__20147\,
            I => \ADC_VDC.n10\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20139\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20134\
        );

    \I__1890\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20134\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__20139\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__20134\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20124\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20119\
        );

    \I__1885\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20119\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__20124\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20119\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__20111\,
            I => \ADC_VDC.n21082\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__20099\,
            I => \ADC_VDC.n21079\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__20096\,
            I => \ADC_VDC.n21977_cascade_\
        );

    \I__1875\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__20090\,
            I => \ADC_VDC.n18482\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20087\,
            I => \bfn_6_6_0_\
        );

    \I__1872\ : InMux
    port map (
            O => \N__20084\,
            I => \ADC_VDC.n19531\
        );

    \I__1871\ : InMux
    port map (
            O => \N__20081\,
            I => \ADC_VDC.n19532\
        );

    \I__1870\ : InMux
    port map (
            O => \N__20078\,
            I => \ADC_VDC.n19533\
        );

    \I__1869\ : InMux
    port map (
            O => \N__20075\,
            I => \ADC_VDC.n19534\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20072\,
            I => \ADC_VDC.n19535\
        );

    \I__1867\ : InMux
    port map (
            O => \N__20069\,
            I => \ADC_VDC.n19536\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20066\,
            I => \ADC_VDC.n19537\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__20063\,
            I => \ADC_IAC.n21068_cascade_\
        );

    \I__1864\ : CEMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__20054\,
            I => \ADC_IAC.n20714\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__1860\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__1856\ : IoSpan4Mux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__20033\,
            I => \IAC_MISO\
        );

    \I__1854\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20024\
        );

    \I__1853\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20024\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__20024\,
            I => cmd_rdadctmp_0_adj_1450
        );

    \I__1851\ : IoInMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__1849\ : Span4Mux_s2_v
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__20008\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__1845\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19999\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__20002\,
            I => \IAC_SCLK\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19999\,
            I => \IAC_SCLK\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__19994\,
            I => \N__19989\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__19993\,
            I => \N__19986\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__19992\,
            I => \N__19983\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19980\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19975\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19975\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19980\,
            I => cmd_rdadctmp_28
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__19975\,
            I => cmd_rdadctmp_28
        );

    \I__1834\ : CEMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__1832\ : Span4Mux_v
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__19958\,
            I => \ADC_IAC.n12\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__19955\,
            I => \n20612_cascade_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19949\,
            I => \ADC_IAC.n20713\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__19946\,
            I => \ADC_IAC.n20783_cascade_\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__19943\,
            I => \ADC_IAC.n20795_cascade_\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__1821\ : Odrv12
    port map (
            O => \N__19931\,
            I => \CLK_DDS.tmp_buf_0\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19924\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19915\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19918\,
            I => bit_cnt_3
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__19915\,
            I => bit_cnt_3
        );

    \I__1814\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19901\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19901\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19901\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19896\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19891\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19891\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__19896\,
            I => bit_cnt_0_adj_1456
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19891\,
            I => bit_cnt_0_adj_1456
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19886\,
            I => \ADC_IAC.n17_cascade_\
        );

    \I__1805\ : IoInMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__1803\ : IoSpan4Mux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1802\ : Span4Mux_s2_v
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__1801\ : Sp12to4
    port map (
            O => \N__19871\,
            I => \N__19867\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__19870\,
            I => \N__19864\
        );

    \I__1799\ : Span12Mux_s11_v
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__1797\ : Odrv12
    port map (
            O => \N__19861\,
            I => \DDS_SCK1\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__19858\,
            I => \DDS_SCK1\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__19853\,
            I => \N__19849\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19844\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19844\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19844\,
            I => cmd_rdadctmp_6_adj_1444
        );

    \I__1791\ : IoInMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1789\ : Span4Mux_s2_v
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__19823\,
            I => \DDS_CS1\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__1782\ : Span12Mux_h
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__1781\ : Span12Mux_v
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__19808\,
            I => \RTD_SDO\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19805\,
            I => \ADC_VDC.n19466\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19802\,
            I => \ADC_VDC.n19467\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19795\
        );

    \I__1776\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19792\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__19795\,
            I => \N__19789\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19792\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__19789\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__1772\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19780\
        );

    \I__1771\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19777\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19774\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__19777\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__19774\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19762\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19759\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__19762\,
            I => \N__19756\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__19759\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__19756\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19747\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19747\,
            I => \N__19741\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__19744\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__19741\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19732\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19729\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19726\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19729\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__19726\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__1751\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19717\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19714\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19711\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__19714\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__1747\ : Odrv12
    port map (
            O => \N__19711\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19699\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19696\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__19699\,
            I => \N__19693\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__19696\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__19693\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19684\
        );

    \I__1739\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19681\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19678\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__19681\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__19678\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__1735\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19670\,
            I => \ADC_VDC.n20\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__19667\,
            I => \ADC_VDC.n19_adj_1412_cascade_\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \ADC_VDC.n18479_cascade_\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19661\,
            I => \ADC_VDC.n19457\
        );

    \I__1730\ : InMux
    port map (
            O => \N__19658\,
            I => \ADC_VDC.n19458\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19655\,
            I => \ADC_VDC.n19459\
        );

    \I__1728\ : InMux
    port map (
            O => \N__19652\,
            I => \ADC_VDC.n19460\
        );

    \I__1727\ : InMux
    port map (
            O => \N__19649\,
            I => \ADC_VDC.n19461\
        );

    \I__1726\ : InMux
    port map (
            O => \N__19646\,
            I => \ADC_VDC.n19462\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19643\,
            I => \ADC_VDC.n19463\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19640\,
            I => \bfn_5_6_0_\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19637\,
            I => \ADC_VDC.n19465\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__19631\,
            I => n20615
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \N__19623\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19620\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__19626\,
            I => \N__19617\
        );

    \I__1717\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19610\
        );

    \I__1716\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19610\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19610\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19605\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19600\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19600\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__19605\,
            I => \N__19595\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19595\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__19589\,
            I => \VAC_DRDY\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__19586\,
            I => \n20615_cascade_\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19576\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19576\
        );

    \I__1703\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19573\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__19576\,
            I => bit_cnt_2
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__19573\,
            I => bit_cnt_2
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19563\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__19567\,
            I => \N__19559\
        );

    \I__1698\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19552\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19552\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19552\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19549\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__19552\,
            I => bit_cnt_1
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__19549\,
            I => bit_cnt_1
        );

    \I__1692\ : SRMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__19535\,
            I => \CLK_DDS.n16766\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19532\,
            I => \bfn_5_5_0_\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \ADC_VAC.n20715_cascade_\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19523\,
            I => \ADC_VAC.n21053\
        );

    \I__1684\ : CEMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19517\,
            I => \ADC_VAC.n20716\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \ADC_VAC.n17_cascade_\
        );

    \I__1681\ : CEMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__19502\,
            I => \ADC_VAC.n12\
        );

    \I__1677\ : CEMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19492\
        );

    \I__1675\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19489\
        );

    \I__1674\ : Span4Mux_h
    port map (
            O => \N__19492\,
            I => \N__19486\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19483\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__19486\,
            I => \ADC_VAC.n12489\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__19483\,
            I => \ADC_VAC.n12489\
        );

    \I__1670\ : IoInMux
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__1668\ : IoSpan4Mux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1667\ : Span4Mux_s2_h
    port map (
            O => \N__19469\,
            I => \N__19465\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__1665\ : Span4Mux_h
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__19459\,
            I => \VAC_SCLK\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19456\,
            I => \VAC_SCLK\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__19451\,
            I => \n14_adj_1606_cascade_\
        );

    \I__1660\ : IoInMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__1658\ : Span4Mux_s2_h
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__19439\,
            I => \N__19435\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__1655\ : Sp12to4
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__1653\ : Odrv12
    port map (
            O => \N__19429\,
            I => \VAC_CS\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__19426\,
            I => \VAC_CS\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19417\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19417\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19414\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19405\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__19405\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__19402\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__19397\,
            I => \ADC_VAC.n21054_cascade_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__19391\,
            I => \ADC_VAC.n16\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1639\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__19370\,
            I => \VAC_MISO\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19361\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19361\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__19361\,
            I => cmd_rdadctmp_0
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19351\
        );

    \I__1628\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__19351\,
            I => cmd_rdadctmp_1
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__19348\,
            I => cmd_rdadctmp_1
        );

    \I__1625\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19337\
        );

    \I__1624\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19337\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__19337\,
            I => cmd_rdadctmp_2
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__19334\,
            I => \N__19330\
        );

    \I__1621\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__1620\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19325\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__19325\,
            I => cmd_rdadctmp_3
        );

    \I__1618\ : SRMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1615\ : Span4Mux_s3_h
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__19310\,
            I => \ADC_VAC.n14822\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19307\,
            I => \ADC_VAC.n19408\
        );

    \I__1612\ : InMux
    port map (
            O => \N__19304\,
            I => \ADC_VAC.n19409\
        );

    \I__1611\ : InMux
    port map (
            O => \N__19301\,
            I => \ADC_VAC.n19410\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19298\,
            I => \ADC_VAC.n19411\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19295\,
            I => \ADC_VAC.n19412\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19292\,
            I => \ADC_VAC.n19413\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19289\,
            I => \ADC_VAC.n19414\
        );

    \I__1606\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19282\
        );

    \I__1605\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__19282\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__19279\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__19274\,
            I => \N__19270\
        );

    \I__1601\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19267\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19264\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__19267\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__19264\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__1597\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19255\
        );

    \I__1596\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19252\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__19255\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19252\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__1593\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19243\
        );

    \I__1592\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19240\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__19243\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__19240\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \N__19231\
        );

    \I__1588\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19228\
        );

    \I__1587\ : InMux
    port map (
            O => \N__19231\,
            I => \N__19225\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__19228\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__19225\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__1584\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19216\
        );

    \I__1583\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19213\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__19216\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__19213\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__1580\ : InMux
    port map (
            O => \N__19208\,
            I => \bfn_2_7_0_\
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1577\ : IoSpan4Mux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__19193\,
            I => \ICE_SYSCLK\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1572\ : IoSpan4Mux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1571\ : Span4Mux_s3_v
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1569\ : Span12Mux_h
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__1568\ : Odrv12
    port map (
            O => \N__19172\,
            I => \ICE_GPMO_2\
        );

    \INVcomm_spi.imiso_83_12208_12209_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12208_12209_resetC_net\,
            I => \N__56995\
        );

    \INVcomm_spi.MISO_48_12202_12203_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12202_12203_setC_net\,
            I => \N__57904\
        );

    \INVcomm_spi.MISO_48_12202_12203_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12202_12203_resetC_net\,
            I => \N__57892\
        );

    \INVcomm_spi.imiso_83_12208_12209_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12208_12209_setC_net\,
            I => \N__56998\
        );

    \INVcomm_spi.bit_cnt_3778__i3C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_3778__i3C_net\,
            I => \N__57036\
        );

    \INVdds0_mclk_304C\ : INV
    port map (
            O => \INVdds0_mclk_304C_net\,
            I => \N__45085\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__57916\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__57899\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__57834\
        );

    \INVADC_VDC.genclk.t_clk_24C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t_clk_24C_net\,
            I => \N__45079\
        );

    \INVdds0_mclkcnt_i7_3783__i0C\ : INV
    port map (
            O => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            I => \N__45082\
        );

    \INVeis_state_i2C\ : INV
    port map (
            O => \INVeis_state_i2C_net\,
            I => \N__57872\
        );

    \INVADC_VDC.genclk.t0on_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i8C_net\,
            I => \N__45078\
        );

    \INVADC_VDC.genclk.t0on_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i0C_net\,
            I => \N__45074\
        );

    \INVADC_VDC.genclk.div_state_i1C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i1C_net\,
            I => \N__45073\
        );

    \INVADC_VDC.genclk.div_state_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i0C_net\,
            I => \N__45072\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__57922\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__57909\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__57894\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__57868\
        );

    \INVeis_end_309C\ : INV
    port map (
            O => \INVeis_end_309C_net\,
            I => \N__57859\
        );

    \INVADC_VDC.genclk.t0off_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i8C_net\,
            I => \N__45071\
        );

    \INVADC_VDC.genclk.t0off_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i0C_net\,
            I => \N__45070\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__57861\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__57851\
        );

    \INViac_raw_buf_vac_raw_buf_merged2WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            I => \N__57932\
        );

    \INViac_raw_buf_vac_raw_buf_merged7WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            I => \N__57983\
        );

    \INViac_raw_buf_vac_raw_buf_merged1WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            I => \N__57857\
        );

    \INViac_raw_buf_vac_raw_buf_merged6WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            I => \N__57981\
        );

    \INViac_raw_buf_vac_raw_buf_merged0WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            I => \N__57838\
        );

    \INViac_raw_buf_vac_raw_buf_merged5WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            I => \N__57978\
        );

    \INViac_raw_buf_vac_raw_buf_merged9WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            I => \N__57847\
        );

    \INViac_raw_buf_vac_raw_buf_merged4WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            I => \N__57969\
        );

    \INViac_raw_buf_vac_raw_buf_merged8WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            I => \N__57828\
        );

    \INViac_raw_buf_vac_raw_buf_merged10WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            I => \N__57878\
        );

    \INViac_raw_buf_vac_raw_buf_merged3WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            I => \N__57955\
        );

    \INViac_raw_buf_vac_raw_buf_merged11WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            I => \N__57906\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19516,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19524,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n19369_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19377,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19361,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19352,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19400,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19391,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_3_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19475\,
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_13_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_5_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19490\,
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19464\,
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_10_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_5_0_\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19429\,
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19437\,
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19445\,
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19453\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \ADC_VAC.bit_cnt_i0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__19208\,
            lcout => \ADC_VAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \ADC_VAC.n19408\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19408\,
            in2 => \_gnd_net_\,
            in3 => \N__19307\,
            lcout => \ADC_VAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19408\,
            carryout => \ADC_VAC.n19409\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19220\,
            in2 => \_gnd_net_\,
            in3 => \N__19304\,
            lcout => \ADC_VAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19409\,
            carryout => \ADC_VAC.n19410\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19247\,
            in2 => \_gnd_net_\,
            in3 => \N__19301\,
            lcout => \ADC_VAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19410\,
            carryout => \ADC_VAC.n19411\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19259\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => \ADC_VAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19411\,
            carryout => \ADC_VAC.n19412\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19234\,
            in2 => \_gnd_net_\,
            in3 => \N__19295\,
            lcout => \ADC_VAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19412\,
            carryout => \ADC_VAC.n19413\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i6_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19273\,
            in2 => \_gnd_net_\,
            in3 => \N__19292\,
            lcout => \ADC_VAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19413\,
            carryout => \ADC_VAC.n19414\,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.bit_cnt_i7_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19421\,
            in2 => \_gnd_net_\,
            in3 => \N__19289\,
            lcout => \ADC_VAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57920\,
            ce => \N__19499\,
            sr => \N__19322\
        );

    \ADC_VAC.i6_4_lut_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__35008\,
            in1 => \N__19285\,
            in2 => \N__19274\,
            in3 => \N__35139\,
            lcout => \ADC_VAC.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19039_4_lut_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19258\,
            in1 => \N__19246\,
            in2 => \N__19235\,
            in3 => \N__19219\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18824_4_lut_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19420\,
            in1 => \N__19409\,
            in2 => \N__19397\,
            in3 => \N__19394\,
            lcout => \ADC_VAC.n21053\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i0_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19366\,
            in1 => \N__34296\,
            in2 => \N__19388\,
            in3 => \N__35215\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i1_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35214\,
            in1 => \N__19367\,
            in2 => \N__34333\,
            in3 => \N__19354\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i4_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35216\,
            in1 => \N__21826\,
            in2 => \N__34332\,
            in3 => \N__19333\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i2_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19342\,
            in1 => \N__34291\,
            in2 => \N__19358\,
            in3 => \N__35217\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i3_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__19343\,
            in1 => \N__34292\,
            in2 => \N__19334\,
            in3 => \N__35218\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57907\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i12409_2_lut_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34938\,
            in2 => \_gnd_net_\,
            in3 => \N__19495\,
            lcout => \ADC_VAC.n14822\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i2_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35166\,
            in2 => \N__34959\,
            in3 => \N__35024\,
            lcout => \DTRIG_N_919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57921\,
            ce => \N__19511\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__35025\,
            in1 => \N__34949\,
            in2 => \_gnd_net_\,
            in3 => \N__35168\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57921\,
            ce => \N__19511\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__34926\,
            in1 => \N__35130\,
            in2 => \N__19626\,
            in3 => \N__32228\,
            lcout => OPEN,
            ltout => \ADC_VAC.n20715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_adj_3_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__35019\,
            in1 => \_gnd_net_\,
            in2 => \N__19529\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC.n20716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i0_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__35165\,
            in1 => \N__35020\,
            in2 => \N__34945\,
            in3 => \N__19526\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57933\,
            ce => \N__19520\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i30_4_lut_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001010001"
        )
    port map (
            in0 => \N__34925\,
            in1 => \N__35018\,
            in2 => \N__19628\,
            in3 => \N__32227\,
            lcout => OPEN,
            ltout => \ADC_VAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19134_2_lut_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__35129\,
            in1 => \_gnd_net_\,
            in2 => \N__19514\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_adj_4_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100010"
        )
    port map (
            in0 => \N__34924\,
            in1 => \N__35128\,
            in2 => \N__19627\,
            in3 => \N__35017\,
            lcout => \ADC_VAC.n12489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.SCLK_35_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011100010"
        )
    port map (
            in0 => \N__34941\,
            in1 => \N__35167\,
            in2 => \N__19468\,
            in3 => \N__35031\,
            lcout => \VAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_140_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__35170\,
            in1 => \N__34940\,
            in2 => \N__19438\,
            in3 => \N__35030\,
            lcout => OPEN,
            ltout => \n14_adj_1606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.CS_37_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__19608\,
            in1 => \N__19634\,
            in2 => \N__19451\,
            in3 => \N__35171\,
            lcout => \VAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_149_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34939\,
            in2 => \_gnd_net_\,
            in3 => \N__35029\,
            lcout => n20615,
            ltout => \n20615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_3_lut_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__19609\,
            in1 => \_gnd_net_\,
            in2 => \N__19586\,
            in3 => \N__35169\,
            lcout => n12534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i2_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23358\,
            lcout => dds_state_2_adj_1452,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i3_3_lut_4_lut_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19581\,
            in1 => \N__23392\,
            in2 => \N__19567\,
            in3 => \N__22543\,
            lcout => n8_adj_1608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i3_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__19583\,
            in1 => \N__19910\,
            in2 => \N__19928\,
            in3 => \N__19566\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57962\,
            ce => \N__23357\,
            sr => \N__19544\
        );

    \CLK_DDS.bit_cnt_i2_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__19909\,
            in1 => \_gnd_net_\,
            in2 => \N__19568\,
            in3 => \N__19582\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57962\,
            ce => \N__23357\,
            sr => \N__19544\
        );

    \CLK_DDS.bit_cnt_i1_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19562\,
            in2 => \_gnd_net_\,
            in3 => \N__19908\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57962\,
            ce => \N__23357\,
            sr => \N__19544\
        );

    \CLK_DDS.i1_3_lut_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__23352\,
            in1 => \N__23421\,
            in2 => \_gnd_net_\,
            in3 => \N__22583\,
            lcout => \CLK_DDS.n16766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.avg_cnt_i0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19720\,
            in2 => \_gnd_net_\,
            in3 => \N__19532\,
            lcout => \ADC_VDC.avg_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \ADC_VDC.n19457\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23815\,
            in2 => \_gnd_net_\,
            in3 => \N__19661\,
            lcout => \ADC_VDC.avg_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19457\,
            carryout => \ADC_VDC.n19458\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23836\,
            in2 => \_gnd_net_\,
            in3 => \N__19658\,
            lcout => \ADC_VDC.avg_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19458\,
            carryout => \ADC_VDC.n19459\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i3_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19765\,
            in2 => \_gnd_net_\,
            in3 => \N__19655\,
            lcout => \ADC_VDC.avg_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19459\,
            carryout => \ADC_VDC.n19460\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19798\,
            in2 => \_gnd_net_\,
            in3 => \N__19652\,
            lcout => \ADC_VDC.avg_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19460\,
            carryout => \ADC_VDC.n19461\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i5_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19750\,
            in2 => \_gnd_net_\,
            in3 => \N__19649\,
            lcout => \ADC_VDC.avg_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19461\,
            carryout => \ADC_VDC.n19462\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i6_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23797\,
            in2 => \_gnd_net_\,
            in3 => \N__19646\,
            lcout => \ADC_VDC.avg_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19462\,
            carryout => \ADC_VDC.n19463\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i7_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19783\,
            in2 => \_gnd_net_\,
            in3 => \N__19643\,
            lcout => \ADC_VDC.avg_cnt_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19463\,
            carryout => \ADC_VDC.n19464\,
            clk => \N__40135\,
            ce => \N__27171\,
            sr => \N__27100\
        );

    \ADC_VDC.avg_cnt_i8_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19702\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \ADC_VDC.avg_cnt_8\,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \ADC_VDC.n19465\,
            clk => \N__40110\,
            ce => \N__27173\,
            sr => \N__27095\
        );

    \ADC_VDC.avg_cnt_i9_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19735\,
            in2 => \_gnd_net_\,
            in3 => \N__19637\,
            lcout => \ADC_VDC.avg_cnt_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19465\,
            carryout => \ADC_VDC.n19466\,
            clk => \N__40110\,
            ce => \N__27173\,
            sr => \N__27095\
        );

    \ADC_VDC.avg_cnt_i10_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19687\,
            in2 => \_gnd_net_\,
            in3 => \N__19805\,
            lcout => \ADC_VDC.avg_cnt_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19466\,
            carryout => \ADC_VDC.n19467\,
            clk => \N__40110\,
            ce => \N__27173\,
            sr => \N__27095\
        );

    \ADC_VDC.avg_cnt_i11_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23854\,
            in2 => \_gnd_net_\,
            in3 => \N__19802\,
            lcout => \ADC_VDC.avg_cnt_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40110\,
            ce => \N__27173\,
            sr => \N__27095\
        );

    \ADC_VDC.i4_4_lut_adj_31_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20971\,
            in1 => \N__20308\,
            in2 => \N__21071\,
            in3 => \N__20170\,
            lcout => \ADC_VDC.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_28_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20258\,
            in2 => \_gnd_net_\,
            in3 => \N__20309\,
            lcout => \ADC_VDC.n6_adj_1410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i8_4_lut_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19799\,
            in1 => \N__19784\,
            in2 => \N__19769\,
            in3 => \N__19751\,
            lcout => \ADC_VDC.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i1_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23319\,
            in1 => \N__23511\,
            in2 => \N__19940\,
            in3 => \N__38398\,
            lcout => \CLK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57879\,
            ce => \N__23177\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7_4_lut_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19736\,
            in1 => \N__19721\,
            in2 => \N__19706\,
            in3 => \N__19688\,
            lcout => OPEN,
            ltout => \ADC_VDC.n19_adj_1412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i11_3_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19673\,
            in2 => \N__19667\,
            in3 => \N__23783\,
            lcout => \ADC_VDC.n18479\,
            ltout => \ADC_VDC.n18479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16053_3_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32859\,
            in2 => \N__19664\,
            in3 => \N__33517\,
            lcout => \ADC_VDC.n18482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i19_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29171\,
            in1 => \N__33372\,
            in2 => \N__23875\,
            in3 => \N__26861\,
            lcout => buf_adcdata_vdc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.CS_28_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__23316\,
            in1 => \N__23488\,
            in2 => \_gnd_net_\,
            in3 => \N__22573\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57908\,
            ce => \N__21755\,
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i11_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__23977\,
            in1 => \N__21545\,
            in2 => \N__21115\,
            in3 => \N__22156\,
            lcout => read_buf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i10_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__22155\,
            in1 => \N__20431\,
            in2 => \N__21560\,
            in3 => \N__23976\,
            lcout => read_buf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.mode_53_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__20321\,
            in1 => \N__21338\,
            in2 => \N__24102\,
            in3 => \N__22397\,
            lcout => \RTD.mode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i12_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__21111\,
            in2 => \N__21561\,
            in3 => \N__20196\,
            lcout => read_buf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24885\,
            in1 => \N__19820\,
            in2 => \N__21559\,
            in3 => \N__22154\,
            lcout => read_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i14_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22159\,
            in1 => \N__23925\,
            in2 => \N__21563\,
            in3 => \N__20524\,
            lcout => read_buf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i15_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__23926\,
            in1 => \N__21546\,
            in2 => \N__21304\,
            in3 => \N__22160\,
            lcout => read_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i13_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22158\,
            in1 => \N__20523\,
            in2 => \N__21562\,
            in3 => \N__20197\,
            lcout => read_buf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23318\,
            in1 => \N__23440\,
            in2 => \N__23537\,
            in3 => \N__27539\,
            lcout => \CLK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57934\,
            ce => \N__23170\,
            sr => \_gnd_net_\
        );

    \i18807_2_lut_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19899\,
            in2 => \_gnd_net_\,
            in3 => \N__19927\,
            lcout => n21227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101000001010"
        )
    port map (
            in0 => \N__19900\,
            in1 => \N__23484\,
            in2 => \N__23353\,
            in3 => \N__22580\,
            lcout => bit_cnt_0_adj_1456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i6_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20459\,
            in1 => \N__52757\,
            in2 => \N__19853\,
            in3 => \N__51983\,
            lcout => cmd_rdadctmp_6_adj_1444,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i30_4_lut_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001010001"
        )
    port map (
            in0 => \N__35856\,
            in1 => \N__35789\,
            in2 => \N__20675\,
            in3 => \N__32213\,
            lcout => OPEN,
            ltout => \ADC_IAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19132_2_lut_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19886\,
            in3 => \N__52756\,
            lcout => \ADC_IAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.SCLK_27_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000110001"
        )
    port map (
            in0 => \N__23317\,
            in1 => \N__23483\,
            in2 => \N__19870\,
            in3 => \N__22582\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i7_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__52758\,
            in2 => \N__25159\,
            in3 => \N__51984\,
            lcout => cmd_rdadctmp_7_adj_1443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_adj_5_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__20670\,
            in1 => \N__35787\,
            in2 => \N__35867\,
            in3 => \N__52707\,
            lcout => \ADC_IAC.n12586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__52708\,
            in1 => \N__35855\,
            in2 => \_gnd_net_\,
            in3 => \N__35786\,
            lcout => \DTRIG_N_919_adj_1451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57963\,
            ce => \N__19970\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i1_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35788\,
            in2 => \N__35868\,
            in3 => \N__52709\,
            lcout => adc_state_1_adj_1417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57963\,
            ce => \N__19970\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_199_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35847\,
            in2 => \_gnd_net_\,
            in3 => \N__35784\,
            lcout => n20612,
            ltout => \n20612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_3_lut_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__20669\,
            in1 => \_gnd_net_\,
            in2 => \N__19955\,
            in3 => \N__52706\,
            lcout => n12663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35851\,
            in2 => \_gnd_net_\,
            in3 => \N__35785\,
            lcout => n20584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_2_lut_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35790\,
            in2 => \_gnd_net_\,
            in3 => \N__19952\,
            lcout => \ADC_IAC.n20714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111101111"
        )
    port map (
            in0 => \N__52720\,
            in1 => \N__35857\,
            in2 => \N__20657\,
            in3 => \N__32226\,
            lcout => \ADC_IAC.n20713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18169_4_lut_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20866\,
            in1 => \N__20545\,
            in2 => \N__20579\,
            in3 => \N__20560\,
            lcout => OPEN,
            ltout => \ADC_IAC.n20783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18181_4_lut_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20836\,
            in1 => \N__20593\,
            in2 => \N__19946\,
            in3 => \N__20818\,
            lcout => OPEN,
            ltout => \ADC_IAC.n20795_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18845_4_lut_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20851\,
            in1 => \N__52721\,
            in2 => \N__19943\,
            in3 => \N__35791\,
            lcout => OPEN,
            ltout => \ADC_IAC.n21068_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i0_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__35792\,
            in1 => \N__52755\,
            in2 => \N__20063\,
            in3 => \N__35858\,
            lcout => adc_state_0_adj_1418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57971\,
            ce => \N__20060\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i1_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52754\,
            in1 => \N__20030\,
            in2 => \N__20774\,
            in3 => \N__52015\,
            lcout => cmd_rdadctmp_1_adj_1449,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i0_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52753\,
            in1 => \N__20029\,
            in2 => \N__20051\,
            in3 => \N__52014\,
            lcout => cmd_rdadctmp_0_adj_1450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.SCLK_35_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__52752\,
            in1 => \N__35869\,
            in2 => \N__20011\,
            in3 => \N__35803\,
            lcout => \IAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i1_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23510\,
            in2 => \_gnd_net_\,
            in3 => \N__22581\,
            lcout => dds_state_1_adj_1453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57979\,
            ce => \N__22492\,
            sr => \N__23359\
        );

    \ADC_VAC.cmd_rdadctmp_i29_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35320\,
            in1 => \N__21909\,
            in2 => \N__19993\,
            in3 => \N__34335\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i28_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35319\,
            in1 => \N__29459\,
            in2 => \N__19992\,
            in3 => \N__34334\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i20_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34653\,
            in1 => \N__35306\,
            in2 => \N__19994\,
            in3 => \N__21942\,
            lcout => buf_adcdata_vac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16066_3_lut_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__33612\,
            in1 => \N__32872\,
            in2 => \_gnd_net_\,
            in3 => \N__33519\,
            lcout => \ADC_VDC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18135_2_lut_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33613\,
            lcout => \ADC_VDC.n20748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i15177_2_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32870\,
            in2 => \_gnd_net_\,
            in3 => \N__33518\,
            lcout => \ADC_VDC.n7_adj_1411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.bit_cnt_3780__i0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20975\,
            in2 => \_gnd_net_\,
            in3 => \N__20087\,
            lcout => \ADC_VDC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \ADC_VDC.n19531\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21070\,
            in2 => \_gnd_net_\,
            in3 => \N__20084\,
            lcout => \ADC_VDC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19531\,
            carryout => \ADC_VDC.n19532\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20314\,
            in2 => \_gnd_net_\,
            in3 => \N__20081\,
            lcout => \ADC_VDC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19532\,
            carryout => \ADC_VDC.n19533\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20267\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \ADC_VDC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19533\,
            carryout => \ADC_VDC.n19534\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i4_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21020\,
            in2 => \_gnd_net_\,
            in3 => \N__20075\,
            lcout => \ADC_VDC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19534\,
            carryout => \ADC_VDC.n19535\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i5_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20171\,
            in2 => \_gnd_net_\,
            in3 => \N__20072\,
            lcout => \ADC_VDC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19535\,
            carryout => \ADC_VDC.n19536\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i6_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20129\,
            in2 => \_gnd_net_\,
            in3 => \N__20069\,
            lcout => \ADC_VDC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19536\,
            carryout => \ADC_VDC.n19537\,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.bit_cnt_3780__i7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20144\,
            in2 => \_gnd_net_\,
            in3 => \N__20066\,
            lcout => \ADC_VDC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40109\,
            ce => \N__33647\,
            sr => \N__21134\
        );

    \ADC_VDC.i18857_4_lut_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__20114\,
            in1 => \N__33521\,
            in2 => \N__21027\,
            in3 => \N__21041\,
            lcout => \ADC_VDC.n21079\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20169\,
            in1 => \N__20142\,
            in2 => \_gnd_net_\,
            in3 => \N__20127\,
            lcout => \ADC_VDC.n20534\,
            ltout => \ADC_VDC.n20534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_3_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111110"
        )
    port map (
            in0 => \N__20972\,
            in1 => \N__21067\,
            in2 => \N__20153\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i5_3_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20150\,
            in1 => \N__20143\,
            in2 => \_gnd_net_\,
            in3 => \N__20128\,
            lcout => \ADC_VDC.n20562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i8_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26621\,
            in1 => \N__30535\,
            in2 => \N__29177\,
            in3 => \N__33346\,
            lcout => buf_adcdata_vdc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i23_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33345\,
            in1 => \N__29173\,
            in2 => \N__22294\,
            in3 => \N__27029\,
            lcout => buf_adcdata_vdc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19094_4_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__21068\,
            in1 => \N__20973\,
            in2 => \N__20268\,
            in3 => \N__20310\,
            lcout => \ADC_VDC.n21082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.n21974_bdd_4_lut_4_lut_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100110000"
        )
    port map (
            in0 => \N__33516\,
            in1 => \N__33349\,
            in2 => \N__20108\,
            in3 => \N__20276\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21977_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33350\,
            in1 => \N__33022\,
            in2 => \N__20096\,
            in3 => \N__20093\,
            lcout => \ADC_VDC.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40111\,
            ce => \N__20213\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__20269\,
            in1 => \N__20315\,
            in2 => \N__21028\,
            in3 => \N__20285\,
            lcout => \ADC_VDC.n10552\,
            ltout => \ADC_VDC.n10552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001001100"
        )
    port map (
            in0 => \N__33348\,
            in1 => \N__32858\,
            in2 => \N__20279\,
            in3 => \N__33515\,
            lcout => \ADC_VDC.n21974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18952_4_lut_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20270\,
            in1 => \N__33011\,
            in2 => \N__21029\,
            in3 => \N__20237\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i37_4_lut_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000110101010"
        )
    port map (
            in0 => \N__33588\,
            in1 => \N__32857\,
            in2 => \N__20228\,
            in3 => \N__33514\,
            lcout => OPEN,
            ltout => \ADC_VDC.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__20225\,
            in1 => \N__33012\,
            in2 => \N__20216\,
            in3 => \N__33347\,
            lcout => \ADC_VDC.n20555\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i6_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__21283\,
            in1 => \N__20490\,
            in2 => \N__20360\,
            in3 => \N__21211\,
            lcout => adress_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i12_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__25408\,
            in1 => \N__24201\,
            in2 => \N__20201\,
            in3 => \N__24473\,
            lcout => \buf_readRTD_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i4_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__20368\,
            in1 => \N__20486\,
            in2 => \N__20183\,
            in3 => \N__21209\,
            lcout => adress_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__21208\,
            in1 => \N__20378\,
            in2 => \N__20491\,
            in3 => \N__20179\,
            lcout => adress_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__20377\,
            in1 => \N__20482\,
            in2 => \N__20414\,
            in3 => \N__21207\,
            lcout => adress_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i5_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__21210\,
            in1 => \N__20369\,
            in2 => \N__20492\,
            in3 => \N__20356\,
            lcout => adress_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.MOSI_59_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__24447\,
            in1 => \N__21238\,
            in2 => \N__21398\,
            in3 => \N__24847\,
            lcout => \RTD_SDI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43815\,
            ce => \N__21347\,
            sr => \N__24514\
        );

    \RTD.i18150_rep_64_2_lut_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24443\,
            in2 => \_gnd_net_\,
            in3 => \N__24843\,
            lcout => \RTD.n22370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19089_3_lut_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__22425\,
            in1 => \N__24845\,
            in2 => \_gnd_net_\,
            in3 => \N__21333\,
            lcout => OPEN,
            ltout => \RTD.n21309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_7_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__24673\,
            in1 => \N__24445\,
            in2 => \N__20324\,
            in3 => \N__22454\,
            lcout => \RTD.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i16303_3_lut_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010101"
        )
    port map (
            in0 => \N__24444\,
            in1 => \_gnd_net_\,
            in2 => \N__22461\,
            in3 => \N__24844\,
            lcout => \RTD.n20762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_11_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24842\,
            in2 => \_gnd_net_\,
            in3 => \N__24664\,
            lcout => \RTD.n20631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i34_4_lut_4_lut_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000111"
        )
    port map (
            in0 => \N__22426\,
            in1 => \N__24846\,
            in2 => \N__25049\,
            in3 => \N__22387\,
            lcout => OPEN,
            ltout => \RTD.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i36_4_lut_4_lut_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000110000"
        )
    port map (
            in0 => \N__22637\,
            in1 => \N__24446\,
            in2 => \N__20435\,
            in3 => \N__24665\,
            lcout => n13181,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i9_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20510\,
            in1 => \N__21524\,
            in2 => \N__20432\,
            in3 => \N__22163\,
            lcout => read_buf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i9_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__24470\,
            in1 => \N__20430\,
            in2 => \N__24235\,
            in3 => \N__27562\,
            lcout => \buf_readRTD_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i1_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__43339\,
            in1 => \N__24222\,
            in2 => \N__20396\,
            in3 => \N__24472\,
            lcout => \buf_readRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__22162\,
            in1 => \N__20394\,
            in2 => \N__21607\,
            in3 => \N__21525\,
            lcout => read_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__38311\,
            in1 => \N__24471\,
            in2 => \N__21587\,
            in3 => \N__24223\,
            lcout => \buf_readRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__20470\,
            in1 => \N__20407\,
            in2 => \N__21227\,
            in3 => \N__21206\,
            lcout => adress_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24893\,
            in1 => \N__21523\,
            in2 => \N__20395\,
            in3 => \N__22161\,
            lcout => read_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12602_2_lut_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24676\,
            in2 => \_gnd_net_\,
            in3 => \N__21376\,
            lcout => \RTD.n15015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i8_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__24468\,
            in1 => \N__25375\,
            in2 => \N__24236\,
            in3 => \N__20506\,
            lcout => \buf_readRTD_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i7_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__21521\,
            in1 => \N__21621\,
            in2 => \N__24259\,
            in3 => \N__22168\,
            lcout => read_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i13_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__25132\,
            in1 => \N__24229\,
            in2 => \N__20531\,
            in3 => \N__24469\,
            lcout => \buf_readRTD_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i8_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22169\,
            in1 => \N__20505\,
            in2 => \N__21628\,
            in3 => \N__21522\,
            lcout => read_buf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i6_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__21464\,
            in2 => \N__24258\,
            in3 => \N__22167\,
            lcout => read_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18141_2_lut_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__25040\,
            in1 => \N__24643\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n20754,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i30_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__51981\,
            in1 => \N__21735\,
            in2 => \N__52916\,
            in3 => \N__21444\,
            lcout => cmd_rdadctmp_30_adj_1420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i29_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20706\,
            in1 => \N__52850\,
            in2 => \N__21448\,
            in3 => \N__51982\,
            lcout => cmd_rdadctmp_29_adj_1421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57935\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i28_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52747\,
            in1 => \N__25297\,
            in2 => \N__20710\,
            in3 => \N__51979\,
            lcout => cmd_rdadctmp_28_adj_1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i5_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__51978\,
            in1 => \N__20458\,
            in2 => \N__20447\,
            in3 => \N__52751\,
            lcout => cmd_rdadctmp_5_adj_1445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i4_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52748\,
            in1 => \N__20443\,
            in2 => \N__20687\,
            in3 => \N__51980\,
            lcout => cmd_rdadctmp_4_adj_1446,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__51977\,
            in1 => \N__20683\,
            in2 => \N__20759\,
            in3 => \N__52750\,
            lcout => cmd_rdadctmp_3_adj_1447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_137_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__52746\,
            in1 => \N__35859\,
            in2 => \N__20611\,
            in3 => \N__35799\,
            lcout => OPEN,
            ltout => \n14_adj_1604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.CS_37_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__20671\,
            in1 => \N__20630\,
            in2 => \N__20624\,
            in3 => \N__52749\,
            lcout => \IAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i12447_2_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35860\,
            in2 => \_gnd_net_\,
            in3 => \N__20797\,
            lcout => \ADC_IAC.n14860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.bit_cnt_i0_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20594\,
            in2 => \_gnd_net_\,
            in3 => \N__20582\,
            lcout => \ADC_IAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \ADC_IAC.n19415\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i1_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20578\,
            in2 => \_gnd_net_\,
            in3 => \N__20564\,
            lcout => \ADC_IAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19415\,
            carryout => \ADC_IAC.n19416\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i2_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20561\,
            in2 => \_gnd_net_\,
            in3 => \N__20549\,
            lcout => \ADC_IAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19416\,
            carryout => \ADC_IAC.n19417\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i3_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20546\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \ADC_IAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19417\,
            carryout => \ADC_IAC.n19418\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i4_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20867\,
            in2 => \_gnd_net_\,
            in3 => \N__20855\,
            lcout => \ADC_IAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19418\,
            carryout => \ADC_IAC.n19419\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i5_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20852\,
            in2 => \_gnd_net_\,
            in3 => \N__20840\,
            lcout => \ADC_IAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19419\,
            carryout => \ADC_IAC.n19420\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i6_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20837\,
            in2 => \_gnd_net_\,
            in3 => \N__20825\,
            lcout => \ADC_IAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19420\,
            carryout => \ADC_IAC.n19421\,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \ADC_IAC.bit_cnt_i7_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20819\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \ADC_IAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57958\,
            ce => \N__20807\,
            sr => \N__20786\
        );

    \CLK_DDS.i19097_4_lut_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100111001100"
        )
    port map (
            in0 => \N__23228\,
            in1 => \N__23489\,
            in2 => \N__23126\,
            in3 => \N__22574\,
            lcout => \CLK_DDS.n12800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i2_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20773\,
            in1 => \N__52819\,
            in2 => \N__20755\,
            in3 => \N__52016\,
            lcout => cmd_rdadctmp_2_adj_1448,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_main.i19670_1_lut_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45097\,
            lcout => \DDS_MCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i20_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53184\,
            in1 => \N__52995\,
            in2 => \N__20720\,
            in3 => \N__40362\,
            lcout => buf_adcdata_iac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__33240\,
            in1 => \N__32896\,
            in2 => \_gnd_net_\,
            in3 => \N__33523\,
            lcout => adc_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40108\,
            ce => \N__20915\,
            sr => \N__20909\
        );

    \ADC_VDC.ADC_DATA_i2_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29131\,
            in1 => \N__33239\,
            in2 => \N__28636\,
            in3 => \N__26315\,
            lcout => buf_adcdata_vdc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i40_3_lut_4_lut_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100100101"
        )
    port map (
            in0 => \N__33492\,
            in1 => \N__32898\,
            in2 => \N__33632\,
            in3 => \N__20947\,
            lcout => OPEN,
            ltout => \ADC_VDC.n19_adj_1413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19163_4_lut_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__33044\,
            in1 => \N__33238\,
            in2 => \N__20918\,
            in3 => \N__20884\,
            lcout => \ADC_VDC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19168_4_lut_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__20894\,
            in1 => \N__33235\,
            in2 => \N__33631\,
            in3 => \N__33043\,
            lcout => \ADC_VDC.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7717_3_lut_4_lut_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111001100"
        )
    port map (
            in0 => \N__20948\,
            in1 => \N__33628\,
            in2 => \N__32906\,
            in3 => \N__33493\,
            lcout => OPEN,
            ltout => \ADC_VDC.n10132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111100"
        )
    port map (
            in0 => \N__20885\,
            in1 => \N__33236\,
            in2 => \N__20897\,
            in3 => \N__33045\,
            lcout => \ADC_VDC.n12823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18137_2_lut_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33621\,
            in2 => \_gnd_net_\,
            in3 => \N__20893\,
            lcout => \ADC_VDC.n20750\,
            ltout => \ADC_VDC.n20750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_32_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111101110"
        )
    port map (
            in0 => \N__20876\,
            in1 => \N__33234\,
            in2 => \N__20870\,
            in3 => \N__33042\,
            lcout => \ADC_VDC.n72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19101_4_lut_4_lut_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110001"
        )
    port map (
            in0 => \N__33476\,
            in1 => \N__32904\,
            in2 => \N__33126\,
            in3 => \N__33283\,
            lcout => OPEN,
            ltout => \ADC_VDC.n11692_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.SCLK_46_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__32905\,
            in1 => \N__21088\,
            in2 => \N__21095\,
            in3 => \N__25820\,
            lcout => \VDC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29110\,
            in1 => \N__33285\,
            in2 => \N__28933\,
            in3 => \N__26348\,
            lcout => buf_adcdata_vdc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21069\,
            in2 => \_gnd_net_\,
            in3 => \N__21040\,
            lcout => OPEN,
            ltout => \ADC_VDC.n11281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_29_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21016\,
            in1 => \N__20990\,
            in2 => \N__20978\,
            in3 => \N__20974\,
            lcout => \ADC_VDC.n15\,
            ltout => \ADC_VDC.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18133_2_lut_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20939\,
            in3 => \N__33475\,
            lcout => OPEN,
            ltout => \ADC_VDC.n20746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_33_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__21146\,
            in1 => \N__32903\,
            in2 => \N__20936\,
            in3 => \N__20933\,
            lcout => \ADC_VDC.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33284\,
            in1 => \N__29111\,
            in2 => \N__23671\,
            in3 => \N__26660\,
            lcout => buf_adcdata_vdc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010010000001100"
        )
    port map (
            in0 => \N__33472\,
            in1 => \N__32988\,
            in2 => \N__33340\,
            in3 => \N__32860\,
            lcout => adc_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40133\,
            ce => \N__20927\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000001000"
        )
    port map (
            in0 => \N__32983\,
            in1 => \N__32845\,
            in2 => \N__33520\,
            in3 => \N__33270\,
            lcout => \ADC_VDC.n13038\,
            ltout => \ADC_VDC.n13038_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i12557_2_lut_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21149\,
            in3 => \N__32985\,
            lcout => \ADC_VDC.n14931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_30_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32984\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33271\,
            lcout => \ADC_VDC.n20659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_36_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32986\,
            lcout => \ADC_VDC.n20392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i15034_2_lut_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33272\,
            in2 => \_gnd_net_\,
            in3 => \N__32846\,
            lcout => OPEN,
            ltout => \ADC_VDC.n17432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_adj_35_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__33471\,
            in1 => \N__32987\,
            in2 => \N__21137\,
            in3 => \N__32768\,
            lcout => \ADC_VDC.n18466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__24140\,
            in1 => \N__24107\,
            in2 => \N__27626\,
            in3 => \N__22316\,
            lcout => \RTD.cfg_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i5_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24110\,
            in1 => \N__24143\,
            in2 => \N__27505\,
            in3 => \N__21182\,
            lcout => \RTD.cfg_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__24142\,
            in1 => \N__24109\,
            in2 => \N__21170\,
            in3 => \N__25205\,
            lcout => \RTD.cfg_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24106\,
            in1 => \N__24139\,
            in2 => \N__25364\,
            in3 => \N__21260\,
            lcout => \RTD.cfg_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i11_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__23902\,
            in1 => \N__24202\,
            in2 => \N__21122\,
            in3 => \N__24436\,
            lcout => \buf_readRTD_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i6_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24108\,
            in1 => \N__24141\,
            in2 => \N__29515\,
            in3 => \N__21272\,
            lcout => \RTD.cfg_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_17_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__24808\,
            in1 => \N__24435\,
            in2 => \N__24680\,
            in3 => \N__25038\,
            lcout => n11730,
            ltout => \n11730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i15_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__24437\,
            in1 => \N__21311\,
            in2 => \N__21287\,
            in3 => \N__22231\,
            lcout => \buf_readRTD_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i7_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__25011\,
            in1 => \N__21284\,
            in2 => \N__24806\,
            in3 => \N__22390\,
            lcout => \RTD.adress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43806\,
            ce => \N__21215\,
            sr => \N__24518\
        );

    \RTD.i1_4_lut_adj_14_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25360\,
            in1 => \N__21271\,
            in2 => \N__29508\,
            in3 => \N__21259\,
            lcout => OPEN,
            ltout => \RTD.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i7_4_lut_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22304\,
            in1 => \N__24914\,
            in2 => \N__21248\,
            in3 => \N__21155\,
            lcout => \RTD.adress_7_N_1340_7\,
            ltout => \RTD.adress_7_N_1340_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24765\,
            in2 => \N__21245\,
            in3 => \N__25009\,
            lcout => \RTD.n20587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__25010\,
            in1 => \N__24799\,
            in2 => \N__21242\,
            in3 => \N__22389\,
            lcout => adress_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43806\,
            ce => \N__21215\,
            sr => \N__24518\
        );

    \RTD.i3_4_lut_adj_13_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25204\,
            in1 => \N__21181\,
            in2 => \N__27506\,
            in3 => \N__21166\,
            lcout => \RTD.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4918_2_lut_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24369\,
            in2 => \_gnd_net_\,
            in3 => \N__25012\,
            lcout => \RTD.n7333\,
            ltout => \RTD.n7333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__24666\,
            in1 => \N__24839\,
            in2 => \N__21353\,
            in3 => \N__22364\,
            lcout => \RTD.n11742\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i30_3_lut_4_lut_3_lut_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24659\,
            in1 => \N__24793\,
            in2 => \_gnd_net_\,
            in3 => \N__25013\,
            lcout => OPEN,
            ltout => \RTD.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i29_4_lut_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__24660\,
            in2 => \N__21350\,
            in3 => \N__22615\,
            lcout => \RTD.n13228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i27_4_lut_4_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110100000010"
        )
    port map (
            in0 => \N__25014\,
            in1 => \N__24841\,
            in2 => \N__24682\,
            in3 => \N__24417\,
            lcout => \RTD.n11734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19144_4_lut_4_lut_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110111111"
        )
    port map (
            in0 => \N__24840\,
            in1 => \N__24371\,
            in2 => \N__24681\,
            in3 => \N__25015\,
            lcout => \RTD.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__24794\,
            in1 => \N__21334\,
            in2 => \N__24683\,
            in3 => \N__22706\,
            lcout => adc_state_1_adj_1483,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43814\,
            ce => \N__22683\,
            sr => \_gnd_net_\
        );

    \RTD.cfg_tmp_i1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__24420\,
            in1 => \N__27615\,
            in2 => \N__24863\,
            in3 => \N__21383\,
            lcout => \RTD.cfg_tmp_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__21317\,
            in1 => \N__24801\,
            in2 => \N__25102\,
            in3 => \N__24427\,
            lcout => \RTD.cfg_tmp_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__24421\,
            in1 => \N__21428\,
            in2 => \N__24864\,
            in3 => \N__25197\,
            lcout => \RTD.cfg_tmp_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i4_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__21422\,
            in1 => \N__24424\,
            in2 => \N__25256\,
            in3 => \N__24849\,
            lcout => \RTD.cfg_tmp_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i5_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__24422\,
            in1 => \N__27501\,
            in2 => \N__24865\,
            in3 => \N__21416\,
            lcout => \RTD.cfg_tmp_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i6_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__21410\,
            in1 => \N__24425\,
            in2 => \N__29516\,
            in3 => \N__24850\,
            lcout => \RTD.cfg_tmp_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__24423\,
            in1 => \N__24065\,
            in2 => \N__24866\,
            in3 => \N__21404\,
            lcout => \RTD.cfg_tmp_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.cfg_tmp_i0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__24800\,
            in2 => \N__25359\,
            in3 => \N__24426\,
            lcout => \RTD.cfg_tmp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43804\,
            ce => \N__21377\,
            sr => \N__21365\
        );

    \RTD.READ_DATA_i4_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__24218\,
            in1 => \N__21478\,
            in2 => \N__38182\,
            in3 => \N__24442\,
            lcout => \buf_readRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__24439\,
            in1 => \N__46891\,
            in2 => \N__21608\,
            in3 => \N__24219\,
            lcout => \buf_readRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__22165\,
            in1 => \N__21477\,
            in2 => \N__21586\,
            in3 => \N__21519\,
            lcout => read_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__24441\,
            in1 => \N__35653\,
            in2 => \N__21629\,
            in3 => \N__24221\,
            lcout => \buf_readRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i3_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__22164\,
            in1 => \N__21606\,
            in2 => \N__21585\,
            in3 => \N__21518\,
            lcout => read_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i5_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__24440\,
            in1 => \N__21463\,
            in2 => \N__43600\,
            in3 => \N__24220\,
            lcout => \buf_readRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_adj_9_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24848\,
            in1 => \N__24584\,
            in2 => \_gnd_net_\,
            in3 => \N__24438\,
            lcout => n1_adj_1601,
            ltout => \n1_adj_1601_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i5_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__21479\,
            in1 => \N__21462\,
            in2 => \N__21467\,
            in3 => \N__22166\,
            lcout => read_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i26_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__22950\,
            in1 => \N__52849\,
            in2 => \N__21667\,
            in3 => \N__52047\,
            lcout => cmd_rdadctmp_26_adj_1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i15_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53127\,
            in1 => \N__52846\,
            in2 => \N__21704\,
            in3 => \N__44949\,
            lcout => buf_adcdata_iac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i21_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53128\,
            in1 => \N__52847\,
            in2 => \N__21449\,
            in3 => \N__22881\,
            lcout => buf_adcdata_iac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i31_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__52046\,
            in1 => \N__21736\,
            in2 => \N__22930\,
            in3 => \N__52854\,
            lcout => cmd_rdadctmp_31_adj_1419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i22_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53129\,
            in1 => \N__52848\,
            in2 => \N__21740\,
            in3 => \N__36795\,
            lcout => buf_adcdata_iac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i27_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52880\,
            in1 => \N__25296\,
            in2 => \N__21668\,
            in3 => \N__52003\,
            lcout => cmd_rdadctmp_27_adj_1423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i16_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53068\,
            in1 => \N__52875\,
            in2 => \N__21686\,
            in3 => \N__22782\,
            lcout => buf_adcdata_iac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.MOSI_31_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23533\,
            in1 => \N__21715\,
            in2 => \_gnd_net_\,
            in3 => \N__23342\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i23_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21699\,
            in1 => \N__52877\,
            in2 => \N__30881\,
            in3 => \N__52004\,
            lcout => cmd_rdadctmp_23_adj_1427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i24_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21700\,
            in1 => \N__52878\,
            in2 => \N__21685\,
            in3 => \N__52005\,
            lcout => cmd_rdadctmp_24_adj_1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i25_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52879\,
            in1 => \N__21681\,
            in2 => \N__22954\,
            in3 => \N__52002\,
            lcout => cmd_rdadctmp_25_adj_1425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i18_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53069\,
            in1 => \N__52876\,
            in2 => \N__27447\,
            in3 => \N__21666\,
            lcout => buf_adcdata_iac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i5_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23333\,
            in1 => \N__23497\,
            in2 => \N__21785\,
            in3 => \N__36302\,
            lcout => \CLK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57947\,
            ce => \N__23145\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i2_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23331\,
            in1 => \N__23496\,
            in2 => \N__21647\,
            in3 => \N__27884\,
            lcout => \CLK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57947\,
            ce => \N__23145\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i3_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__23495\,
            in1 => \N__23334\,
            in2 => \N__21803\,
            in3 => \N__27656\,
            lcout => \CLK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57947\,
            ce => \N__23145\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i4_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__23332\,
            in1 => \N__25745\,
            in2 => \N__21794\,
            in3 => \N__23498\,
            lcout => \CLK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57947\,
            ce => \N__23145\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i6_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__23494\,
            in2 => \N__31286\,
            in3 => \N__23326\,
            lcout => \CLK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57959\,
            ce => \N__23144\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i7_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23325\,
            in1 => \N__23499\,
            in2 => \N__21770\,
            in3 => \N__44588\,
            lcout => \CLK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57959\,
            ce => \N__23144\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i8_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__21761\,
            in1 => \N__23327\,
            in2 => \N__23513\,
            in3 => \N__25592\,
            lcout => \CLK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57959\,
            ce => \N__23144\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.i23_4_lut_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000010011"
        )
    port map (
            in0 => \N__22575\,
            in1 => \N__23323\,
            in2 => \N__23121\,
            in3 => \N__23490\,
            lcout => \CLK_DDS.n9_adj_1395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19153_4_lut_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__23324\,
            in1 => \N__22576\,
            in2 => \N__23512\,
            in3 => \N__23114\,
            lcout => \CLK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i12_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__25968\,
            in1 => \N__34454\,
            in2 => \N__28835\,
            in3 => \N__35305\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i4_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__25972\,
            in1 => \N__34658\,
            in2 => \N__35423\,
            in3 => \N__21886\,
            lcout => buf_adcdata_vac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i4_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53185\,
            in1 => \N__52996\,
            in2 => \N__28763\,
            in3 => \N__21862\,
            lcout => buf_adcdata_iac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_5_i22_3_lut_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21983\,
            in1 => \N__25861\,
            in2 => \_gnd_net_\,
            in3 => \N__49056\,
            lcout => n22_adj_1632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_4_i19_3_lut_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22043\,
            in1 => \N__21885\,
            in2 => \_gnd_net_\,
            in3 => \N__56358\,
            lcout => OPEN,
            ltout => \n19_adj_1636_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_4_i22_3_lut_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49057\,
            in1 => \_gnd_net_\,
            in2 => \N__21872\,
            in3 => \N__21861\,
            lcout => OPEN,
            ltout => \n22_adj_1637_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_4_i30_3_lut_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21848\,
            in2 => \N__21836\,
            in3 => \N__48669\,
            lcout => n30_adj_1638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i16_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35368\,
            in1 => \N__21994\,
            in2 => \N__30576\,
            in3 => \N__34337\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i5_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__34338\,
            in1 => \N__35372\,
            in2 => \N__21815\,
            in3 => \N__21833\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i21_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35366\,
            in1 => \N__34657\,
            in2 => \N__21923\,
            in3 => \N__25470\,
            lcout => buf_adcdata_vac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i7_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34656\,
            in1 => \N__35371\,
            in2 => \N__21998\,
            in3 => \N__23650\,
            lcout => buf_adcdata_vac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i6_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35369\,
            in1 => \N__21814\,
            in2 => \N__25921\,
            in3 => \N__34339\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i6_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34655\,
            in1 => \N__35370\,
            in2 => \N__23590\,
            in3 => \N__23695\,
            lcout => buf_adcdata_vac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i15_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35367\,
            in1 => \N__21993\,
            in2 => \N__23696\,
            in3 => \N__34336\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_5_i19_3_lut_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21969\,
            in1 => \N__56295\,
            in2 => \_gnd_net_\,
            in3 => \N__22058\,
            lcout => n19_adj_1631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i5_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35361\,
            in1 => \N__34661\,
            in2 => \N__25952\,
            in3 => \N__21973\,
            lcout => buf_adcdata_vac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i23_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34660\,
            in1 => \N__35364\,
            in2 => \N__22073\,
            in3 => \N__22263\,
            lcout => buf_adcdata_vac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__33237\,
            in2 => \N__33124\,
            in3 => \N__33491\,
            lcout => n13109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22202_bdd_4_lut_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__25397\,
            in1 => \N__21943\,
            in2 => \N__22028\,
            in3 => \N__48419\,
            lcout => n22205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i22_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34659\,
            in1 => \N__35363\,
            in2 => \N__31965\,
            in3 => \N__22087\,
            lcout => buf_adcdata_vac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i30_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35362\,
            in1 => \N__21922\,
            in2 => \N__22088\,
            in3 => \N__34439\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i31_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__34440\,
            in1 => \N__22086\,
            in2 => \N__22072\,
            in3 => \N__35365\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i5_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33294\,
            in1 => \N__22054\,
            in2 => \N__29162\,
            in3 => \N__26744\,
            lcout => buf_adcdata_vdc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__30484\,
            in1 => \N__33295\,
            in2 => \N__26552\,
            in3 => \N__29124\,
            lcout => buf_adcdata_vdc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i4_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__22039\,
            in2 => \N__29161\,
            in3 => \N__26786\,
            lcout => buf_adcdata_vdc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i17_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__43978\,
            in1 => \N__29125\,
            in2 => \N__26903\,
            in3 => \N__33296\,
            lcout => buf_adcdata_vdc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i20_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__22021\,
            in2 => \N__29159\,
            in3 => \N__27239\,
            lcout => buf_adcdata_vdc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i6_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__23557\,
            in1 => \N__33298\,
            in2 => \N__26705\,
            in3 => \N__29127\,
            lcout => buf_adcdata_vdc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33292\,
            in1 => \N__28510\,
            in2 => \N__29160\,
            in3 => \N__26825\,
            lcout => buf_adcdata_vdc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i21_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__25435\,
            in1 => \N__29126\,
            in2 => \N__27218\,
            in3 => \N__33297\,
            lcout => buf_adcdata_vdc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110110"
        )
    port map (
            in0 => \N__33344\,
            in1 => \N__33086\,
            in2 => \N__33614\,
            in3 => \N__33477\,
            lcout => \ADC_VDC.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40136\,
            ce => \N__22010\,
            sr => \_gnd_net_\
        );

    \i15243_2_lut_3_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__37981\,
            in1 => \_gnd_net_\,
            in2 => \N__54172\,
            in3 => \N__52436\,
            lcout => n14_adj_1579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15253_2_lut_3_lut_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__52437\,
            in1 => \N__54145\,
            in2 => \_gnd_net_\,
            in3 => \N__43149\,
            lcout => n14_adj_1570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15255_2_lut_3_lut_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__52435\,
            in1 => \N__54141\,
            in2 => \_gnd_net_\,
            in3 => \N__44291\,
            lcout => n14_adj_1572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15256_2_lut_3_lut_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__42971\,
            in1 => \_gnd_net_\,
            in2 => \N__54173\,
            in3 => \N__52439\,
            lcout => n14_adj_1573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15257_2_lut_3_lut_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52438\,
            in1 => \N__45545\,
            in2 => \_gnd_net_\,
            in3 => \N__54149\,
            lcout => n14_adj_1574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.SCLK_51_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100100011100"
        )
    port map (
            in0 => \N__24805\,
            in1 => \N__24434\,
            in2 => \N__24679\,
            in3 => \N__25034\,
            lcout => \RTD_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43816\,
            ce => \N__22181\,
            sr => \_gnd_net_\
        );

    \RTD.i19171_4_lut_4_lut_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011110111000"
        )
    port map (
            in0 => \N__24802\,
            in1 => \N__24431\,
            in2 => \N__24677\,
            in3 => \N__25031\,
            lcout => \RTD.n11756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_4_lut_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000110"
        )
    port map (
            in0 => \N__25030\,
            in1 => \N__24644\,
            in2 => \N__24467\,
            in3 => \N__24803\,
            lcout => \RTD.n15081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_16_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010110001"
        )
    port map (
            in0 => \N__24804\,
            in1 => \N__24433\,
            in2 => \N__24678\,
            in3 => \N__25033\,
            lcout => n13309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19100_3_lut_3_lut_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__24648\,
            in1 => \N__24432\,
            in2 => \_gnd_net_\,
            in3 => \N__25032\,
            lcout => \RTD.n11703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_15_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22430\,
            in2 => \_gnd_net_\,
            in3 => \N__22388\,
            lcout => \RTD.n16669\,
            ltout => \RTD.n16669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.CS_52_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001101110111"
        )
    port map (
            in0 => \N__25039\,
            in1 => \N__24658\,
            in2 => \N__22358\,
            in3 => \N__24797\,
            lcout => \RTD_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43780\,
            ce => \N__22334\,
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__24022\,
            in1 => \N__24063\,
            in2 => \N__27622\,
            in3 => \N__22315\,
            lcout => \RTD.n12_adj_1397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16108_3_lut_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__22264\,
            in2 => \_gnd_net_\,
            in3 => \N__56248\,
            lcout => OPEN,
            ltout => \n19_adj_1526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19474_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__22220\,
            in1 => \N__48398\,
            in2 => \N__22244\,
            in3 => \N__49054\,
            lcout => OPEN,
            ltout => \n22076_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22076_bdd_4_lut_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49055\,
            in1 => \N__24491\,
            in2 => \N__22241\,
            in3 => \N__22805\,
            lcout => n22079,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i20_3_lut_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56247\,
            in1 => \N__22238\,
            in2 => \_gnd_net_\,
            in3 => \N__24062\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__22652\,
            in1 => \N__22214\,
            in2 => \N__24675\,
            in3 => \N__22727\,
            lcout => \RTD.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43740\,
            ce => \N__22684\,
            sr => \_gnd_net_\
        );

    \RTD.i19088_2_lut_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__25017\,
            in1 => \N__33845\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \RTD.n21323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i45_4_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000100010"
        )
    port map (
            in0 => \N__24411\,
            in1 => \N__22632\,
            in2 => \N__22655\,
            in3 => \N__31703\,
            lcout => \RTD.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19023_4_lut_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__22643\,
            in1 => \N__24636\,
            in2 => \N__22468\,
            in3 => \N__22721\,
            lcout => OPEN,
            ltout => \RTD.n21325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__24413\,
            in1 => \N__22633\,
            in2 => \N__22646\,
            in3 => \N__24635\,
            lcout => adc_state_2_adj_1482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43740\,
            ce => \N__22684\,
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_12_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__25018\,
            in1 => \_gnd_net_\,
            in2 => \N__24807\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4948_2_lut_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24769\,
            in2 => \_gnd_net_\,
            in3 => \N__25016\,
            lcout => \RTD.n1\,
            ltout => \RTD.n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_4_lut_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000110000000"
        )
    port map (
            in0 => \N__24634\,
            in1 => \N__24412\,
            in2 => \N__22619\,
            in3 => \N__22616\,
            lcout => \RTD.n13192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001100000011"
        )
    port map (
            in0 => \N__22604\,
            in1 => \N__22532\,
            in2 => \N__23360\,
            in3 => \N__22595\,
            lcout => dds_state_0_adj_1454,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57881\,
            ce => \N__22493\,
            sr => \_gnd_net_\
        );

    \RTD.i18725_4_lut_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24409\,
            in1 => \N__25019\,
            in2 => \N__22469\,
            in3 => \N__22720\,
            lcout => OPEN,
            ltout => \RTD.n21276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19037_3_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24795\,
            in2 => \N__22730\,
            in3 => \N__24928\,
            lcout => \RTD.n21275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33840\,
            in2 => \_gnd_net_\,
            in3 => \N__31701\,
            lcout => \RTD.adc_state_3_N_1368_1\,
            ltout => \RTD.adc_state_3_N_1368_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100111101110"
        )
    port map (
            in0 => \N__24410\,
            in1 => \N__24798\,
            in2 => \N__22709\,
            in3 => \N__25020\,
            lcout => \RTD.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__24466\,
            in1 => \N__24591\,
            in2 => \N__22700\,
            in3 => \N__24929\,
            lcout => adc_state_3_adj_1481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43758\,
            ce => \N__22685\,
            sr => \_gnd_net_\
        );

    \i15266_2_lut_3_lut_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__41499\,
            in1 => \N__54171\,
            in2 => \_gnd_net_\,
            in3 => \N__52433\,
            lcout => n14_adj_1545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_3_i16_3_lut_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28287\,
            in1 => \_gnd_net_\,
            in2 => \N__27655\,
            in3 => \N__56286\,
            lcout => OPEN,
            ltout => \n16_adj_1512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18264_3_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__53230\,
            in1 => \_gnd_net_\,
            in2 => \N__22658\,
            in3 => \N__48374\,
            lcout => n20878,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18225_3_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23011\,
            in1 => \N__56287\,
            in2 => \_gnd_net_\,
            in3 => \N__32345\,
            lcout => n20839,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_218_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__53591\,
            in1 => \N__48503\,
            in2 => \_gnd_net_\,
            in3 => \N__31882\,
            lcout => n20670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i3_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49871\,
            in1 => \N__28288\,
            in2 => \N__37985\,
            in3 => \N__38967\,
            lcout => buf_dds0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i17_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53130\,
            in1 => \N__52845\,
            in2 => \N__22955\,
            in3 => \N__25545\,
            lcout => buf_adcdata_iac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41370\,
            in1 => \N__46059\,
            in2 => \N__49915\,
            in3 => \N__22819\,
            lcout => \VAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i6_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__22906\,
            in1 => \N__41371\,
            in2 => \N__46421\,
            in3 => \N__49875\,
            lcout => \VAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i23_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__52844\,
            in1 => \N__53131\,
            in2 => \N__22931\,
            in3 => \N__22849\,
            lcout => buf_adcdata_iac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19469_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__22905\,
            in1 => \N__48373\,
            in2 => \N__22882\,
            in3 => \N__56246\,
            lcout => n22100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14314_3_lut_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56245\,
            in1 => \N__22848\,
            in2 => \_gnd_net_\,
            in3 => \N__22818\,
            lcout => n17_adj_1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19444_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__22743\,
            in1 => \N__48375\,
            in2 => \N__22783\,
            in3 => \N__56304\,
            lcout => n22040,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22744\,
            in1 => \N__44477\,
            in2 => \_gnd_net_\,
            in3 => \N__41388\,
            lcout => \IAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22100_bdd_4_lut_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48376\,
            in1 => \N__28117\,
            in2 => \N__23033\,
            in3 => \N__30994\,
            lcout => n22103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i5_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__30942\,
            in1 => \N__44430\,
            in2 => \N__49925\,
            in3 => \N__46406\,
            lcout => \AMPV_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i7_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28979\,
            in1 => \N__49910\,
            in2 => \N__46067\,
            in3 => \N__24047\,
            lcout => \buf_cfgRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i2_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49909\,
            in1 => \N__44429\,
            in2 => \N__43005\,
            in3 => \N__23007\,
            lcout => \SELIRNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_4_i16_3_lut_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56305\,
            in1 => \N__25740\,
            in2 => \_gnd_net_\,
            in3 => \N__28414\,
            lcout => n16_adj_1508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i10_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23335\,
            in1 => \N__23506\,
            in2 => \N__23186\,
            in3 => \N__25798\,
            lcout => \CLK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i11_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__23503\,
            in1 => \N__23339\,
            in2 => \N__22988\,
            in3 => \N__40483\,
            lcout => \CLK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i12_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23336\,
            in1 => \N__23507\,
            in2 => \N__22979\,
            in3 => \N__40293\,
            lcout => \CLK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i13_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23337\,
            in1 => \N__23508\,
            in2 => \N__22970\,
            in3 => \N__30995\,
            lcout => \CLK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i14_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__23340\,
            in2 => \N__36964\,
            in3 => \N__22961\,
            lcout => \CLK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i15_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__23338\,
            in1 => \N__23509\,
            in2 => \N__23546\,
            in3 => \N__25280\,
            lcout => tmp_buf_15_adj_1455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i9_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__23341\,
            in2 => \N__23195\,
            in3 => \N__25609\,
            lcout => \CLK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57937\,
            ce => \N__23169\,
            sr => \_gnd_net_\
        );

    \trig_dds1_315_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__49904\,
            in1 => \N__54981\,
            in2 => \N__23125\,
            in3 => \N__34796\,
            lcout => trig_dds1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_219_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010000"
        )
    port map (
            in0 => \N__34829\,
            in1 => \N__49900\,
            in2 => \N__54983\,
            in3 => \N__36587\,
            lcout => n12411,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i13_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49918\,
            in1 => \N__28116\,
            in2 => \N__46420\,
            in3 => \N__38957\,
            lcout => buf_dds0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i4_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__38955\,
            in1 => \N__51183\,
            in2 => \N__49923\,
            in3 => \N__28413\,
            lcout => buf_dds0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48360\,
            in1 => \N__56360\,
            in2 => \N__34834\,
            in3 => \N__49100\,
            lcout => n20673,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i9_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__38956\,
            in1 => \N__49919\,
            in2 => \N__45576\,
            in3 => \N__28030\,
            lcout => buf_dds0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ICE_GPMO_1_I_0_3_lut_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31373\,
            in1 => \N__23093\,
            in2 => \_gnd_net_\,
            in3 => \N__35720\,
            lcout => \IAC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i14_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35417\,
            in1 => \N__23686\,
            in2 => \N__25948\,
            in3 => \N__34455\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i7_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53199\,
            in1 => \N__52994\,
            in2 => \N__23717\,
            in3 => \N__23623\,
            lcout => buf_adcdata_iac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_7_i19_3_lut_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23675\,
            in1 => \N__23646\,
            in2 => \_gnd_net_\,
            in3 => \N__56359\,
            lcout => OPEN,
            ltout => \n19_adj_1625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_7_i22_3_lut_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23622\,
            in2 => \N__23609\,
            in3 => \N__49116\,
            lcout => OPEN,
            ltout => \n22_adj_1626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_7_i30_3_lut_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__48723\,
            in1 => \N__23606\,
            in2 => \N__23594\,
            in3 => \_gnd_net_\,
            lcout => n30_adj_1627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34654\,
            in1 => \N__35418\,
            in2 => \N__33957\,
            in3 => \N__26970\,
            lcout => buf_adcdata_vac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i13_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52951\,
            in1 => \N__25878\,
            in2 => \N__28762\,
            in3 => \N__52073\,
            lcout => cmd_rdadctmp_13_adj_1437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i6_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__53198\,
            in1 => \N__23767\,
            in2 => \N__52997\,
            in3 => \N__23731\,
            lcout => buf_adcdata_iac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_6_i19_3_lut_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23583\,
            in1 => \N__23564\,
            in2 => \_gnd_net_\,
            in3 => \N__56361\,
            lcout => OPEN,
            ltout => \n19_adj_1628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_6_i22_3_lut_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23766\,
            in2 => \N__23750\,
            in3 => \N__49117\,
            lcout => OPEN,
            ltout => \n22_adj_1629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_6_i30_3_lut_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23747\,
            in2 => \N__23735\,
            in3 => \N__48668\,
            lcout => n30_adj_1630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i14_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__52071\,
            in1 => \N__23727\,
            in2 => \N__25885\,
            in3 => \N__52953\,
            lcout => cmd_rdadctmp_14_adj_1436,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i15_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52952\,
            in1 => \N__23709\,
            in2 => \N__23732\,
            in3 => \N__52074\,
            lcout => cmd_rdadctmp_15_adj_1435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i16_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__52072\,
            in1 => \N__52105\,
            in2 => \N__23716\,
            in3 => \N__52954\,
            lcout => cmd_rdadctmp_16_adj_1434,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__26242\,
            in2 => \N__26180\,
            in3 => \N__26151\,
            lcout => cmd_rdadctmp_1_adj_1478,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i7_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26001\,
            in1 => \N__26520\,
            in2 => \N__26277\,
            in3 => \N__33121\,
            lcout => cmd_rdadctmp_7_adj_1472,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i6_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__33117\,
            in1 => \N__26002\,
            in2 => \N__26036\,
            in3 => \N__26246\,
            lcout => cmd_rdadctmp_6_adj_1473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__26241\,
            in1 => \N__26175\,
            in2 => \N__33629\,
            in3 => \N__33119\,
            lcout => cmd_rdadctmp_0_adj_1479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i9_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33118\,
            in1 => \N__26492\,
            in2 => \N__26459\,
            in3 => \N__26250\,
            lcout => cmd_rdadctmp_9_adj_1470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26031\,
            in1 => \N__26065\,
            in2 => \N__26276\,
            in3 => \N__33120\,
            lcout => cmd_rdadctmp_5_adj_1474,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i12_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33339\,
            in1 => \N__35614\,
            in2 => \N__29163\,
            in3 => \N__26933\,
            lcout => buf_adcdata_vdc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__33109\,
            in1 => \N__26392\,
            in2 => \N__26426\,
            in3 => \N__26232\,
            lcout => cmd_rdadctmp_11_adj_1468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26391\,
            in1 => \N__26364\,
            in2 => \N__26274\,
            in3 => \N__33113\,
            lcout => cmd_rdadctmp_12_adj_1467,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_27_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__33108\,
            in1 => \N__32902\,
            in2 => \N__33358\,
            in3 => \N__33473\,
            lcout => n12875,
            ltout => \n12875_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26330\,
            in1 => \N__26842\,
            in2 => \N__23774\,
            in3 => \N__33114\,
            lcout => cmd_rdadctmp_14_adj_1465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__33110\,
            in1 => \N__26236\,
            in2 => \N__26371\,
            in3 => \N__26329\,
            lcout => cmd_rdadctmp_13_adj_1466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i19_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26637\,
            in1 => \N__26680\,
            in2 => \N__26275\,
            in3 => \N__33115\,
            lcout => cmd_rdadctmp_19_adj_1460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33111\,
            in1 => \N__26638\,
            in2 => \N__26603\,
            in3 => \N__26240\,
            lcout => cmd_rdadctmp_20_adj_1459,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i10_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26421\,
            in1 => \N__26454\,
            in2 => \N__26273\,
            in3 => \N__33112\,
            lcout => cmd_rdadctmp_10_adj_1469,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i18_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__26879\,
            in1 => \N__29150\,
            in2 => \N__23956\,
            in3 => \N__33338\,
            lcout => buf_adcdata_vdc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i11_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33337\,
            in1 => \N__38248\,
            in2 => \N__29172\,
            in3 => \N__26948\,
            lcout => buf_adcdata_vdc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22214_bdd_4_lut_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__48340\,
            in1 => \N__29428\,
            in2 => \N__23882\,
            in3 => \N__23891\,
            lcout => n20828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i15_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26802\,
            in1 => \N__26843\,
            in2 => \N__26278\,
            in3 => \N__33083\,
            lcout => cmd_rdadctmp_15_adj_1464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i17_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__33082\,
            in1 => \N__26721\,
            in2 => \N__26768\,
            in3 => \N__26255\,
            lcout => cmd_rdadctmp_17_adj_1462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26487\,
            in1 => \N__26525\,
            in2 => \N__26280\,
            in3 => \N__33085\,
            lcout => cmd_rdadctmp_8_adj_1471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i16_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33081\,
            in1 => \N__26803\,
            in2 => \N__26767\,
            in3 => \N__26254\,
            lcout => cmd_rdadctmp_16_adj_1463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i18_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26722\,
            in1 => \N__26679\,
            in2 => \N__26279\,
            in3 => \N__33084\,
            lcout => cmd_rdadctmp_18_adj_1461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i9_4_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__23858\,
            in1 => \N__23840\,
            in2 => \N__23822\,
            in3 => \N__23801\,
            lcout => \ADC_VDC.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18888_3_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__27022\,
            in1 => \N__33354\,
            in2 => \_gnd_net_\,
            in3 => \N__24011\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i34_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33123\,
            in1 => \N__27002\,
            in2 => \N__24002\,
            in3 => \N__32867\,
            lcout => cmd_rdadcbuf_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40088\,
            ce => \N__23999\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010101010"
        )
    port map (
            in0 => \N__33122\,
            in1 => \N__32866\,
            in2 => \N__33371\,
            in3 => \N__33474\,
            lcout => \ADC_VDC.n13050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i10_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24418\,
            in1 => \N__24233\,
            in2 => \N__23990\,
            in3 => \N__25120\,
            lcout => \buf_readRTD_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12112_2_lut_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__54106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54846\,
            lcout => n14522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18219_3_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23963\,
            in1 => \N__29029\,
            in2 => \_gnd_net_\,
            in3 => \N__56250\,
            lcout => OPEN,
            ltout => \n20833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19484_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__25058\,
            in1 => \N__48309\,
            in2 => \N__23939\,
            in3 => \N__49059\,
            lcout => n22118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i14_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__24419\,
            in1 => \N__24234\,
            in2 => \N__23936\,
            in3 => \N__28885\,
            lcout => \buf_readRTD_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19562_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56249\,
            in1 => \N__25196\,
            in2 => \N__23912\,
            in3 => \N__48308\,
            lcout => n22214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_4_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25103\,
            in1 => \N__24484\,
            in2 => \N__25255\,
            in3 => \N__24904\,
            lcout => \RTD.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24103\,
            in1 => \N__24125\,
            in2 => \N__25095\,
            in3 => \N__24905\,
            lcout => \RTD.cfg_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__24449\,
            in1 => \N__24892\,
            in2 => \N__41251\,
            in3 => \N__24227\,
            lcout => \buf_readRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_4_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__24796\,
            in1 => \N__24448\,
            in2 => \N__25048\,
            in3 => \N__24674\,
            lcout => \RTD.n14717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i16_3_lut_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25276\,
            in1 => \N__28064\,
            in2 => \_gnd_net_\,
            in3 => \N__56180\,
            lcout => n16_adj_1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24104\,
            in1 => \N__24126\,
            in2 => \N__25248\,
            in3 => \N__24485\,
            lcout => \RTD.cfg_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i6_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__24450\,
            in1 => \N__38044\,
            in2 => \N__24266\,
            in3 => \N__24228\,
            lcout => \buf_readRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__24127\,
            in1 => \N__24105\,
            in2 => \N__24026\,
            in3 => \N__24064\,
            lcout => \RTD.cfg_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__40802\,
            in1 => \N__32053\,
            in2 => \N__48620\,
            in3 => \N__32099\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__44307\,
            in1 => \N__29001\,
            in2 => \N__49917\,
            in3 => \N__25187\,
            lcout => \buf_cfgRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__52089\,
            in1 => \N__25163\,
            in2 => \N__29394\,
            in3 => \N__52911\,
            lcout => cmd_rdadctmp_8_adj_1442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__25085\,
            in1 => \N__29000\,
            in2 => \N__49916\,
            in3 => \N__43009\,
            lcout => \buf_cfgRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19542_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56263\,
            in1 => \N__27473\,
            in2 => \N__25142\,
            in3 => \N__48299\,
            lcout => n22184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18220_3_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25121\,
            in1 => \N__25084\,
            in2 => \_gnd_net_\,
            in3 => \N__56264\,
            lcout => n20834,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_adj_19_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__33844\,
            in1 => \N__25047\,
            in2 => \_gnd_net_\,
            in3 => \N__31702\,
            lcout => \RTD.n20656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_216_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__46609\,
            in1 => \N__54922\,
            in2 => \N__49895\,
            in3 => \N__34830\,
            lcout => n12397,
            ltout => \n12397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__43161\,
            in1 => \N__49839\,
            in2 => \N__24917\,
            in3 => \N__36843\,
            lcout => \VAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_251_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__27672\,
            in1 => \N__27255\,
            in2 => \_gnd_net_\,
            in3 => \N__27270\,
            lcout => n20646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22184_bdd_4_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__48344\,
            in1 => \N__25483\,
            in2 => \N__25448\,
            in3 => \N__25424\,
            lcout => n20849,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19552_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25228\,
            in1 => \N__48342\,
            in2 => \N__25418\,
            in3 => \N__56281\,
            lcout => n22202,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49838\,
            in1 => \N__28996\,
            in2 => \N__45581\,
            in3 => \N__27596\,
            lcout => \buf_cfgRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19395_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25340\,
            in1 => \N__48343\,
            in2 => \N__25385\,
            in3 => \N__56282\,
            lcout => n22016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44467\,
            in1 => \N__28994\,
            in2 => \_gnd_net_\,
            in3 => \N__25332\,
            lcout => \buf_cfgRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i19_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53166\,
            in1 => \N__52915\,
            in2 => \N__25313\,
            in3 => \N__40893\,
            lcout => buf_adcdata_iac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i15_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__25275\,
            in1 => \N__38574\,
            in2 => \N__46066\,
            in3 => \N__38479\,
            lcout => buf_dds1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49921\,
            in1 => \N__28995\,
            in2 => \N__44174\,
            in3 => \N__25229\,
            lcout => \buf_cfgRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__27399\,
            in1 => \N__41375\,
            in2 => \N__43010\,
            in3 => \N__49922\,
            lcout => \IAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22106_bdd_4_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__25571\,
            in1 => \N__25505\,
            in2 => \N__25565\,
            in3 => \N__48538\,
            lcout => n22109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19405_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__48297\,
            in1 => \N__27703\,
            in2 => \N__25546\,
            in3 => \N__56301\,
            lcout => n22022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18262_4_lut_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__48298\,
            in1 => \N__25523\,
            in2 => \N__32153\,
            in3 => \N__56302\,
            lcout => OPEN,
            ltout => \n20876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19479_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25499\,
            in1 => \N__48574\,
            in2 => \N__25508\,
            in3 => \N__49058\,
            lcout => n22106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i12_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__40294\,
            in1 => \N__38573\,
            in2 => \N__44168\,
            in3 => \N__38472\,
            lcout => buf_dds1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_1_i16_3_lut_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56303\,
            in1 => \N__38399\,
            in2 => \_gnd_net_\,
            in3 => \N__28339\,
            lcout => n16_adj_1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18261_4_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__48296\,
            in1 => \N__56300\,
            in2 => \N__30923\,
            in3 => \N__47555\,
            lcout => n20875,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__27845\,
            in1 => \N__54949\,
            in2 => \N__49823\,
            in3 => \N__27836\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22022_bdd_4_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__25608\,
            in1 => \N__25493\,
            in2 => \N__48424\,
            in3 => \N__28023\,
            lcout => n22025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__25744\,
            in1 => \N__38562\,
            in2 => \N__51188\,
            in3 => \N__38455\,
            lcout => buf_dds1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6394_3_lut_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41498\,
            in1 => \N__27920\,
            in2 => \_gnd_net_\,
            in3 => \N__41749\,
            lcout => n8_adj_1555,
            ltout => \n8_adj_1555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_8_i15_4_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49734\,
            in1 => \N__54948\,
            in2 => \N__25724\,
            in3 => \N__27898\,
            lcout => \data_index_9_N_216_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__27899\,
            in1 => \N__49735\,
            in2 => \N__54977\,
            in3 => \N__25625\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22040_bdd_4_lut_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__25587\,
            in1 => \N__25619\,
            in2 => \N__28372\,
            in3 => \N__48377\,
            lcout => n22043,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i10_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__25802\,
            in1 => \N__38557\,
            in2 => \N__43004\,
            in3 => \N__38448\,
            lcout => buf_dds1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i9_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__38450\,
            in1 => \N__25610\,
            in2 => \N__45577\,
            in3 => \N__38563\,
            lcout => buf_dds1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i8_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__25591\,
            in1 => \N__38558\,
            in2 => \N__41510\,
            in3 => \N__38449\,
            lcout => buf_dds1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49899\,
            in1 => \N__38932\,
            in2 => \N__45467\,
            in3 => \N__28335\,
            lcout => buf_dds0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i15_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__28060\,
            in1 => \N__49897\,
            in2 => \N__46058\,
            in3 => \N__38935\,
            lcout => buf_dds0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_213_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__49896\,
            in1 => \N__25781\,
            in2 => \_gnd_net_\,
            in3 => \N__54963\,
            lcout => n12383,
            ltout => \n12383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i8_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__41506\,
            in1 => \N__49898\,
            in2 => \N__25805\,
            in3 => \N__28368\,
            lcout => buf_dds0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18210_3_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25797\,
            in1 => \N__28143\,
            in2 => \_gnd_net_\,
            in3 => \N__56339\,
            lcout => n20824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i2_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__38933\,
            in1 => \N__49914\,
            in2 => \N__47150\,
            in3 => \N__28440\,
            lcout => buf_dds0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i10_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__28144\,
            in1 => \N__49908\,
            in2 => \N__43003\,
            in3 => \N__38934\,
            lcout => buf_dds0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_253_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__51589\,
            in1 => \N__25780\,
            in2 => \N__49924\,
            in3 => \N__54964\,
            lcout => OPEN,
            ltout => \n11412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds0_314_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__54965\,
            in1 => \N__44789\,
            in2 => \N__25769\,
            in3 => \N__49920\,
            lcout => trig_dds0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_I_0_1_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36359\,
            lcout => \AC_ADC_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i8_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__25901\,
            in1 => \N__34424\,
            in2 => \N__26971\,
            in3 => \N__35421\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i13_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__25944\,
            in1 => \N__34456\,
            in2 => \N__25979\,
            in3 => \N__35420\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i7_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35419\,
            in1 => \N__25900\,
            in2 => \N__34460\,
            in3 => \N__25922\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i2_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53206\,
            in1 => \N__52993\,
            in2 => \N__28676\,
            in3 => \N__28585\,
            lcout => buf_adcdata_iac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i5_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__52992\,
            in1 => \N__53207\,
            in2 => \N__25889\,
            in3 => \N__25860\,
            lcout => buf_adcdata_iac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_5_i30_3_lut_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__25841\,
            in1 => \N__25829\,
            in2 => \N__48741\,
            in3 => \_gnd_net_\,
            lcout => n30_adj_1634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i2_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33100\,
            in1 => \N__26121\,
            in2 => \N__26291\,
            in3 => \N__26152\,
            lcout => cmd_rdadctmp_2_adj_1477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i22_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__26569\,
            in1 => \N__31782\,
            in2 => \N__33127\,
            in3 => \N__26284\,
            lcout => cmd_rdadctmp_22_adj_1457,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19104_2_lut_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33301\,
            in2 => \_gnd_net_\,
            in3 => \N__33098\,
            lcout => \ADC_VDC.n21718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i21_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__33099\,
            in1 => \N__26568\,
            in2 => \N__26290\,
            in3 => \N__26602\,
            lcout => cmd_rdadctmp_21_adj_1458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i4_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__26289\,
            in1 => \N__33101\,
            in2 => \N__26096\,
            in3 => \N__26064\,
            lcout => cmd_rdadctmp_4_adj_1475,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i3_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__26122\,
            in1 => \N__26091\,
            in2 => \N__33128\,
            in3 => \N__26288\,
            lcout => cmd_rdadctmp_3_adj_1476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26159\,
            in2 => \N__26179\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.cmd_rdadcbuf_0\,
            ltout => OPEN,
            carryin => \bfn_10_5_0_\,
            carryout => \ADC_VDC.n19422\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26132\,
            in2 => \N__26153\,
            in3 => \N__26126\,
            lcout => \ADC_VDC.cmd_rdadcbuf_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19422\,
            carryout => \ADC_VDC.n19423\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26105\,
            in2 => \N__26123\,
            in3 => \N__26099\,
            lcout => \ADC_VDC.cmd_rdadcbuf_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19423\,
            carryout => \ADC_VDC.n19424\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i3_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26075\,
            in2 => \N__26095\,
            in3 => \N__26069\,
            lcout => \ADC_VDC.cmd_rdadcbuf_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19424\,
            carryout => \ADC_VDC.n19425\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i4_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26045\,
            in2 => \N__26066\,
            in3 => \N__26039\,
            lcout => \ADC_VDC.cmd_rdadcbuf_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19425\,
            carryout => \ADC_VDC.n19426\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26012\,
            in2 => \N__26035\,
            in3 => \N__26006\,
            lcout => \ADC_VDC.cmd_rdadcbuf_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19426\,
            carryout => \ADC_VDC.n19427\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i6_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25985\,
            in2 => \N__26003\,
            in3 => \N__26528\,
            lcout => \ADC_VDC.cmd_rdadcbuf_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19427\,
            carryout => \ADC_VDC.n19428\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i7_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26501\,
            in2 => \N__26524\,
            in3 => \N__26495\,
            lcout => \ADC_VDC.cmd_rdadcbuf_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19428\,
            carryout => \ADC_VDC.n19429\,
            clk => \N__40034\,
            ce => \N__27190\,
            sr => \N__27107\
        );

    \ADC_VDC.cmd_rdadcbuf_i8_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26468\,
            in2 => \N__26491\,
            in3 => \N__26462\,
            lcout => \ADC_VDC.cmd_rdadcbuf_8\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \ADC_VDC.n19430\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i9_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26435\,
            in2 => \N__26458\,
            in3 => \N__26429\,
            lcout => \ADC_VDC.cmd_rdadcbuf_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19430\,
            carryout => \ADC_VDC.n19431\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i10_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26402\,
            in2 => \N__26425\,
            in3 => \N__26396\,
            lcout => \ADC_VDC.cmd_rdadcbuf_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19431\,
            carryout => \ADC_VDC.n19432\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i11_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29200\,
            in2 => \N__26393\,
            in3 => \N__26375\,
            lcout => cmd_rdadcbuf_11,
            ltout => OPEN,
            carryin => \ADC_VDC.n19432\,
            carryout => \ADC_VDC.n19433\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i12_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26344\,
            in2 => \N__26372\,
            in3 => \N__26333\,
            lcout => cmd_rdadcbuf_12,
            ltout => OPEN,
            carryin => \ADC_VDC.n19433\,
            carryout => \ADC_VDC.n19434\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i13_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26328\,
            in2 => \N__26311\,
            in3 => \N__26294\,
            lcout => cmd_rdadcbuf_13,
            ltout => OPEN,
            carryin => \ADC_VDC.n19434\,
            carryout => \ADC_VDC.n19435\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i14_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26841\,
            in2 => \N__26824\,
            in3 => \N__26807\,
            lcout => cmd_rdadcbuf_14,
            ltout => OPEN,
            carryin => \ADC_VDC.n19435\,
            carryout => \ADC_VDC.n19436\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i15_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26782\,
            in2 => \N__26804\,
            in3 => \N__26771\,
            lcout => cmd_rdadcbuf_15,
            ltout => OPEN,
            carryin => \ADC_VDC.n19436\,
            carryout => \ADC_VDC.n19437\,
            clk => \N__40049\,
            ce => \N__27183\,
            sr => \N__27106\
        );

    \ADC_VDC.cmd_rdadcbuf_i16_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26737\,
            in2 => \N__26766\,
            in3 => \N__26726\,
            lcout => cmd_rdadcbuf_16,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \ADC_VDC.n19438\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i17_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26695\,
            in2 => \N__26723\,
            in3 => \N__26684\,
            lcout => cmd_rdadcbuf_17,
            ltout => OPEN,
            carryin => \ADC_VDC.n19438\,
            carryout => \ADC_VDC.n19439\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i18_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26653\,
            in2 => \N__26681\,
            in3 => \N__26642\,
            lcout => cmd_rdadcbuf_18,
            ltout => OPEN,
            carryin => \ADC_VDC.n19439\,
            carryout => \ADC_VDC.n19440\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i19_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26617\,
            in2 => \N__26639\,
            in3 => \N__26606\,
            lcout => cmd_rdadcbuf_19,
            ltout => OPEN,
            carryin => \ADC_VDC.n19440\,
            carryout => \ADC_VDC.n19441\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i20_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29044\,
            in2 => \N__26601\,
            in3 => \N__26576\,
            lcout => cmd_rdadcbuf_20,
            ltout => OPEN,
            carryin => \ADC_VDC.n19441\,
            carryout => \ADC_VDC.n19442\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i21_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26542\,
            in2 => \N__26573\,
            in3 => \N__26531\,
            lcout => cmd_rdadcbuf_21,
            ltout => OPEN,
            carryin => \ADC_VDC.n19442\,
            carryout => \ADC_VDC.n19443\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i22_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26947\,
            in2 => \N__31789\,
            in3 => \N__26936\,
            lcout => cmd_rdadcbuf_22,
            ltout => OPEN,
            carryin => \ADC_VDC.n19443\,
            carryout => \ADC_VDC.n19444\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i23_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26929\,
            in2 => \N__31751\,
            in3 => \N__26918\,
            lcout => cmd_rdadcbuf_23,
            ltout => OPEN,
            carryin => \ADC_VDC.n19444\,
            carryout => \ADC_VDC.n19445\,
            clk => \N__40117\,
            ce => \N__27159\,
            sr => \N__27105\
        );

    \ADC_VDC.cmd_rdadcbuf_i24_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28846\,
            in2 => \_gnd_net_\,
            in3 => \N__26915\,
            lcout => cmd_rdadcbuf_24,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \ADC_VDC.n19446\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i25_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28858\,
            in2 => \_gnd_net_\,
            in3 => \N__26912\,
            lcout => cmd_rdadcbuf_25,
            ltout => OPEN,
            carryin => \ADC_VDC.n19446\,
            carryout => \ADC_VDC.n19447\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i26_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28870\,
            in2 => \_gnd_net_\,
            in3 => \N__26909\,
            lcout => cmd_rdadcbuf_26,
            ltout => OPEN,
            carryin => \ADC_VDC.n19447\,
            carryout => \ADC_VDC.n19448\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i27_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29215\,
            in2 => \_gnd_net_\,
            in3 => \N__26906\,
            lcout => cmd_rdadcbuf_27,
            ltout => OPEN,
            carryin => \ADC_VDC.n19448\,
            carryout => \ADC_VDC.n19449\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i28_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26893\,
            in2 => \_gnd_net_\,
            in3 => \N__26882\,
            lcout => cmd_rdadcbuf_28,
            ltout => OPEN,
            carryin => \ADC_VDC.n19449\,
            carryout => \ADC_VDC.n19450\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i29_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26875\,
            in2 => \_gnd_net_\,
            in3 => \N__26864\,
            lcout => cmd_rdadcbuf_29,
            ltout => OPEN,
            carryin => \ADC_VDC.n19450\,
            carryout => \ADC_VDC.n19451\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i30_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26857\,
            in2 => \_gnd_net_\,
            in3 => \N__26846\,
            lcout => cmd_rdadcbuf_30,
            ltout => OPEN,
            carryin => \ADC_VDC.n19451\,
            carryout => \ADC_VDC.n19452\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i31_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27232\,
            in2 => \_gnd_net_\,
            in3 => \N__27221\,
            lcout => cmd_rdadcbuf_31,
            ltout => OPEN,
            carryin => \ADC_VDC.n19452\,
            carryout => \ADC_VDC.n19453\,
            clk => \N__40116\,
            ce => \N__27172\,
            sr => \N__27099\
        );

    \ADC_VDC.cmd_rdadcbuf_i32_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27208\,
            in2 => \_gnd_net_\,
            in3 => \N__27197\,
            lcout => cmd_rdadcbuf_32,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \ADC_VDC.n19454\,
            clk => \N__40119\,
            ce => \N__27191\,
            sr => \N__27104\
        );

    \ADC_VDC.cmd_rdadcbuf_i33_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29188\,
            in2 => \_gnd_net_\,
            in3 => \N__27194\,
            lcout => cmd_rdadcbuf_33,
            ltout => OPEN,
            carryin => \ADC_VDC.n19454\,
            carryout => \ADC_VDC.n19455\,
            clk => \N__40119\,
            ce => \N__27191\,
            sr => \N__27104\
        );

    \ADC_VDC.add_23_36_lut_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27021\,
            in2 => \_gnd_net_\,
            in3 => \N__27005\,
            lcout => \ADC_VDC.cmd_rdadcbuf_35_N_1139_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_376_i9_2_lut_3_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__48171\,
            in1 => \N__56182\,
            in2 => \_gnd_net_\,
            in3 => \N__48952\,
            lcout => n9_adj_1416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i10_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__34761\,
            in1 => \N__34380\,
            in2 => \N__28531\,
            in3 => \N__35345\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22118_bdd_4_lut_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48953\,
            in1 => \N__27380\,
            in2 => \N__26996\,
            in3 => \N__26978\,
            lcout => n22121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_194_i9_2_lut_3_lut_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__48170\,
            in1 => \N__56181\,
            in2 => \_gnd_net_\,
            in3 => \N__48951\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i9_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__26972\,
            in1 => \N__34382\,
            in2 => \N__34765\,
            in3 => \N__35347\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i5_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49828\,
            in1 => \N__29006\,
            in2 => \N__27483\,
            in3 => \N__46405\,
            lcout => \buf_cfgRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i25_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__29239\,
            in1 => \N__34381\,
            in2 => \N__34482\,
            in3 => \N__35346\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18211_3_lut_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56166\,
            in1 => \N__27451\,
            in2 => \_gnd_net_\,
            in3 => \N__27403\,
            lcout => n20825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i14_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__38964\,
            in1 => \N__43153\,
            in2 => \N__49825\,
            in3 => \N__36909\,
            lcout => buf_dds0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_0_i16_3_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__56167\,
            in1 => \_gnd_net_\,
            in2 => \N__27538\,
            in3 => \N__31189\,
            lcout => n16_adj_1488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_0_i15_4_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54923\,
            in1 => \N__31013\,
            in2 => \N__49824\,
            in3 => \N__30896\,
            lcout => \data_index_9_N_216_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15049_2_lut_3_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__27673\,
            in1 => \N__27256\,
            in2 => \_gnd_net_\,
            in3 => \N__27271\,
            lcout => \comm_state_3_N_436_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__32045\,
            in1 => \N__32101\,
            in2 => \N__51059\,
            in3 => \N__27272\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__40247\,
            in1 => \N__27257\,
            in2 => \N__32116\,
            in3 => \N__32046\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__45544\,
            in1 => \N__49749\,
            in2 => \N__41382\,
            in3 => \N__27693\,
            lcout => \IAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__32122\,
            in1 => \N__32054\,
            in2 => \N__40661\,
            in3 => \N__27674\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i3_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__27648\,
            in1 => \N__38578\,
            in2 => \N__47841\,
            in3 => \N__54946\,
            lcout => buf_dds1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__27595\,
            in1 => \N__48341\,
            in2 => \N__27572\,
            in3 => \N__56159\,
            lcout => n22226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_210_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__27551\,
            in1 => \N__54945\,
            in2 => \N__49826\,
            in3 => \N__46571\,
            lcout => n11931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53175\,
            in1 => \N__52989\,
            in2 => \N__29398\,
            in3 => \N__34051\,
            lcout => buf_adcdata_iac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i14_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__38571\,
            in1 => \N__43168\,
            in2 => \N__36954\,
            in3 => \N__38471\,
            lcout => buf_dds1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__38470\,
            in1 => \N__41163\,
            in2 => \N__27537\,
            in3 => \N__38572\,
            lcout => buf_dds1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_240_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__53568\,
            in1 => \N__48537\,
            in2 => \_gnd_net_\,
            in3 => \N__31880\,
            lcout => n20663,
            ltout => \n20663_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__53995\,
            in1 => \N__52378\,
            in2 => \N__27731\,
            in3 => \N__36582\,
            lcout => n10614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_243_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__56144\,
            in1 => \N__48536\,
            in2 => \_gnd_net_\,
            in3 => \N__31881\,
            lcout => n11354,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15263_2_lut_3_lut_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__53997\,
            in1 => \_gnd_net_\,
            in2 => \N__46028\,
            in3 => \N__52380\,
            lcout => n14_adj_1544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49754\,
            in1 => \N__31188\,
            in2 => \N__41168\,
            in3 => \N__38965\,
            lcout => buf_dds0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15302_2_lut_3_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53996\,
            in1 => \N__41162\,
            in2 => \_gnd_net_\,
            in3 => \N__52379\,
            lcout => n14_adj_1533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_2_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__31031\,
            in1 => \N__31029\,
            in2 => \N__39136\,
            in3 => \N__27728\,
            lcout => n7_adj_1531,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => n19384,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_3_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38606\,
            in1 => \N__38605\,
            in2 => \N__39140\,
            in3 => \N__27725\,
            lcout => n7_adj_1566,
            ltout => OPEN,
            carryin => n19384,
            carryout => n19385,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_4_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36182\,
            in1 => \N__36181\,
            in2 => \N__39137\,
            in3 => \N__27722\,
            lcout => n7_adj_1564,
            ltout => OPEN,
            carryin => n19385,
            carryout => n19386,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_5_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36047\,
            in1 => \N__36046\,
            in2 => \N__39141\,
            in3 => \N__27719\,
            lcout => n7_adj_1562,
            ltout => OPEN,
            carryin => n19386,
            carryout => n19387,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_6_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38768\,
            in1 => \N__38767\,
            in2 => \N__39138\,
            in3 => \N__27716\,
            lcout => n7_adj_1560,
            ltout => OPEN,
            carryin => n19387,
            carryout => n19388,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_7_lut_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__31051\,
            in1 => \N__31050\,
            in2 => \N__39142\,
            in3 => \N__27929\,
            lcout => n17409,
            ltout => OPEN,
            carryin => n19388,
            carryout => n19389,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_8_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41963\,
            in1 => \N__41962\,
            in2 => \N__39139\,
            in3 => \N__27926\,
            lcout => n7_adj_1558,
            ltout => OPEN,
            carryin => n19389,
            carryout => n19390,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_9_lut_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27862\,
            in1 => \N__27861\,
            in2 => \N__39143\,
            in3 => \N__27923\,
            lcout => n7_adj_1556,
            ltout => OPEN,
            carryin => n19390,
            carryout => n19391,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_10_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27919\,
            in1 => \N__27912\,
            in2 => \N__39153\,
            in3 => \N__27890\,
            lcout => n7_adj_1554,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => n19392,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_131_11_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__27985\,
            in1 => \N__27986\,
            in2 => \N__39158\,
            in3 => \N__27887\,
            lcout => n7_adj_1552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_2_i16_3_lut_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27879\,
            in1 => \N__28442\,
            in2 => \_gnd_net_\,
            in3 => \N__56309\,
            lcout => n16_adj_1515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i2_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__27883\,
            in1 => \N__38559\,
            in2 => \N__47143\,
            in3 => \N__38451\,
            lcout => buf_dds1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6404_3_lut_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47672\,
            in1 => \N__27863\,
            in2 => \_gnd_net_\,
            in3 => \N__41709\,
            lcout => n8_adj_1557,
            ltout => \n8_adj_1557_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_7_i15_4_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49830\,
            in1 => \N__54953\,
            in2 => \N__27839\,
            in3 => \N__27835\,
            lcout => \data_index_9_N_216_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6384_3_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45521\,
            in1 => \N__27984\,
            in2 => \_gnd_net_\,
            in3 => \N__41708\,
            lcout => n8_adj_1553,
            ltout => \n8_adj_1553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i9_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49831\,
            in1 => \N__54954\,
            in2 => \N__27989\,
            in3 => \N__28255\,
            lcout => data_index_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_response_312_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001001010010"
        )
    port map (
            in0 => \N__54976\,
            in1 => \N__52389\,
            in2 => \N__54140\,
            in3 => \N__53590\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57926\,
            ce => \N__27944\,
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_297_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000110010"
        )
    port map (
            in0 => \N__53589\,
            in1 => \N__52416\,
            in2 => \N__51590\,
            in3 => \N__54975\,
            lcout => n11401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_227_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__51585\,
            in1 => \N__39482\,
            in2 => \_gnd_net_\,
            in3 => \N__54971\,
            lcout => n11866,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18158_2_lut_3_lut_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54090\,
            in1 => \N__52387\,
            in2 => \_gnd_net_\,
            in3 => \N__53587\,
            lcout => OPEN,
            ltout => \n20772_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_183_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__51584\,
            in1 => \N__54973\,
            in2 => \N__27935\,
            in3 => \N__34795\,
            lcout => n11835,
            ltout => \n11835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_69_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101111"
        )
    port map (
            in0 => \N__54974\,
            in1 => \N__54005\,
            in2 => \N__27932\,
            in3 => \N__52388\,
            lcout => n16763,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_282_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__53588\,
            in1 => \N__54091\,
            in2 => \_gnd_net_\,
            in3 => \N__54972\,
            lcout => n11377,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i14_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__50306\,
            in1 => \N__50138\,
            in2 => \N__36925\,
            in3 => \N__28097\,
            lcout => \SIG_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i11_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50133\,
            in1 => \N__50303\,
            in2 => \N__28130\,
            in3 => \N__40457\,
            lcout => \SIG_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i10_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50302\,
            in1 => \N__50132\,
            in2 => \N__28007\,
            in3 => \N__28145\,
            lcout => \SIG_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i13_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50137\,
            in1 => \N__50305\,
            in2 => \N__28085\,
            in3 => \N__28121\,
            lcout => \SIG_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i6_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50308\,
            in1 => \N__50140\,
            in2 => \N__28451\,
            in3 => \N__31301\,
            lcout => \SIG_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i12_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__40333\,
            in1 => \N__28091\,
            in2 => \N__50157\,
            in3 => \N__50304\,
            lcout => \SIG_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i15_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50307\,
            in1 => \N__50139\,
            in2 => \N__28073\,
            in3 => \N__28056\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i9_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50141\,
            in1 => \N__50309\,
            in2 => \N__28352\,
            in3 => \N__28034\,
            lcout => \SIG_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57939\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i7_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50184\,
            in1 => \N__50300\,
            in2 => \N__27998\,
            in3 => \N__44567\,
            lcout => \SIG_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i5_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__50299\,
            in1 => \N__50183\,
            in2 => \N__28391\,
            in3 => \N__36548\,
            lcout => \SIG_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i2_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50180\,
            in1 => \N__50296\,
            in2 => \N__28316\,
            in3 => \N__28441\,
            lcout => \SIG_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__50298\,
            in1 => \N__50182\,
            in2 => \N__28421\,
            in3 => \N__28271\,
            lcout => \SIG_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i8_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50185\,
            in1 => \N__50301\,
            in2 => \N__28382\,
            in3 => \N__28373\,
            lcout => \SIG_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i1_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__50295\,
            in1 => \N__28340\,
            in2 => \N__31409\,
            in3 => \N__50179\,
            lcout => \SIG_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i3_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50181\,
            in1 => \N__50297\,
            in2 => \N__28307\,
            in3 => \N__28298\,
            lcout => \SIG_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57950\,
            ce => \N__31390\,
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_9_i15_4_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54982\,
            in1 => \N__28265\,
            in2 => \N__49829\,
            in3 => \N__28256\,
            lcout => \data_index_9_N_216_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i2_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34652\,
            in1 => \N__35410\,
            in2 => \N__28541\,
            in3 => \N__28606\,
            lcout => buf_adcdata_vac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31324\,
            in1 => \N__31429\,
            in2 => \N__31472\,
            in3 => \N__31447\,
            lcout => \ADC_VDC.genclk.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_2_i19_3_lut_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28643\,
            in1 => \N__28605\,
            in2 => \_gnd_net_\,
            in3 => \N__56341\,
            lcout => OPEN,
            ltout => \n19_adj_1646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_2_i22_3_lut_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28581\,
            in2 => \N__28565\,
            in3 => \N__49098\,
            lcout => OPEN,
            ltout => \n22_adj_1647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_2_i30_3_lut_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28562\,
            in2 => \N__28544\,
            in3 => \N__48719\,
            lcout => n30_adj_1648,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i11_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35409\,
            in1 => \N__28537\,
            in2 => \N__28824\,
            in3 => \N__34453\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19102_2_lut_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33677\,
            in2 => \_gnd_net_\,
            in3 => \N__40171\,
            lcout => \ADC_VDC.genclk.n11751\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_3_i19_3_lut_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28514\,
            in1 => \N__28794\,
            in2 => \_gnd_net_\,
            in3 => \N__56291\,
            lcout => OPEN,
            ltout => \n19_adj_1642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_3_i22_3_lut_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28464\,
            in2 => \N__28493\,
            in3 => \N__49052\,
            lcout => OPEN,
            ltout => \n22_adj_1643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_3_i30_3_lut_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28490\,
            in2 => \N__28475\,
            in3 => \N__48681\,
            lcout => n30_adj_1644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53200\,
            in1 => \N__52999\,
            in2 => \N__28781\,
            in3 => \N__28465\,
            lcout => buf_adcdata_iac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i3_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34621\,
            in1 => \N__35412\,
            in2 => \N__28834\,
            in3 => \N__28795\,
            lcout => buf_adcdata_vac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i11_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__52077\,
            in1 => \N__28669\,
            in2 => \N__28780\,
            in3 => \N__53000\,
            lcout => cmd_rdadctmp_11_adj_1439,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i12_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52998\,
            in1 => \N__28776\,
            in2 => \N__28755\,
            in3 => \N__52078\,
            lcout => cmd_rdadctmp_12_adj_1438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i17_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35411\,
            in1 => \N__30580\,
            in2 => \N__30430\,
            in3 => \N__34452\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i7_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51406\,
            in1 => \N__28724\,
            in2 => \_gnd_net_\,
            in3 => \N__54138\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57816\,
            ce => \N__31493\,
            sr => \N__31673\
        );

    \comm_buf_5__i6_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54136\,
            in1 => \N__40245\,
            in2 => \_gnd_net_\,
            in3 => \N__28706\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57816\,
            ce => \N__31493\,
            sr => \N__31673\
        );

    \comm_buf_5__i5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51055\,
            in1 => \N__28691\,
            in2 => \_gnd_net_\,
            in3 => \N__54137\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57816\,
            ce => \N__31493\,
            sr => \N__31673\
        );

    \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__29365\,
            in1 => \N__52958\,
            in2 => \N__28668\,
            in3 => \N__52090\,
            lcout => cmd_rdadctmp_10_adj_1440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i36_4_lut_4_lut_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011110100"
        )
    port map (
            in0 => \N__56252\,
            in1 => \N__48195\,
            in2 => \N__48718\,
            in3 => \N__48997\,
            lcout => OPEN,
            ltout => \n30_adj_1480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_96_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__48998\,
            in1 => \N__48266\,
            in2 => \N__28940\,
            in3 => \N__45187\,
            lcout => \comm_state_3_N_420_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_1_i19_3_lut_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56253\,
            in1 => \N__28937\,
            in2 => \_gnd_net_\,
            in3 => \N__34741\,
            lcout => OPEN,
            ltout => \n19_adj_1491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_1_i22_3_lut_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__48999\,
            in1 => \_gnd_net_\,
            in2 => \N__28916\,
            in3 => \N__28905\,
            lcout => n22_adj_1489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__28906\,
            in1 => \N__53183\,
            in2 => \N__29369\,
            in3 => \N__52959\,
            lcout => buf_adcdata_iac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19528_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__48194\,
            in1 => \N__29495\,
            in2 => \N__28892\,
            in3 => \N__56251\,
            lcout => n22160,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i15_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29165\,
            in1 => \N__33366\,
            in2 => \N__29341\,
            in3 => \N__28871\,
            lcout => buf_adcdata_vdc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i14_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33363\,
            in1 => \N__29169\,
            in2 => \N__38101\,
            in3 => \N__28859\,
            lcout => buf_adcdata_vdc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i13_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29164\,
            in1 => \N__33365\,
            in2 => \N__46666\,
            in3 => \N__28847\,
            lcout => buf_adcdata_vdc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_37_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011100000"
        )
    port map (
            in0 => \N__33125\,
            in1 => \N__32868\,
            in2 => \N__33373\,
            in3 => \N__33522\,
            lcout => \ADC_VDC.n12915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i16_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29166\,
            in1 => \N__33367\,
            in2 => \N__29278\,
            in3 => \N__29216\,
            lcout => buf_adcdata_vdc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33362\,
            in1 => \N__29168\,
            in2 => \N__33982\,
            in3 => \N__29204\,
            lcout => buf_adcdata_vdc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i22_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__29167\,
            in1 => \N__29189\,
            in2 => \N__33374\,
            in3 => \N__31924\,
            lcout => buf_adcdata_vdc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i9_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__33364\,
            in1 => \N__29170\,
            in2 => \N__30850\,
            in3 => \N__29045\,
            lcout => buf_adcdata_vdc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_166_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__52432\,
            in1 => \N__54902\,
            in2 => \N__51569\,
            in3 => \N__40496\,
            lcout => n11918,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i18_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34583\,
            in1 => \N__35392\,
            in2 => \N__34244\,
            in3 => \N__29028\,
            lcout => buf_adcdata_vac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__43303\,
            in1 => \N__54903\,
            in2 => \N__47248\,
            in3 => \N__51319\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i6_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__51320\,
            in1 => \N__43201\,
            in2 => \N__54961\,
            in3 => \N__40246\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i27_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35391\,
            in1 => \N__34240\,
            in2 => \N__29451\,
            in3 => \N__34432\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__29005\,
            in1 => \N__49628\,
            in2 => \N__43175\,
            in3 => \N__29488\,
            lcout => \buf_cfgRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i19_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35390\,
            in1 => \N__34584\,
            in2 => \N__29452\,
            in3 => \N__29421\,
            lcout => buf_adcdata_vac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__29399\,
            in1 => \N__52991\,
            in2 => \N__29364\,
            in3 => \N__52094\,
            lcout => cmd_rdadctmp_9_adj_1441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i15_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__29311\,
            in1 => \N__34595\,
            in2 => \N__29261\,
            in3 => \N__35342\,
            lcout => buf_adcdata_vac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_7_i19_3_lut_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29345\,
            in1 => \N__29310\,
            in2 => \_gnd_net_\,
            in3 => \N__55943\,
            lcout => n19_adj_1502,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22016_bdd_4_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__30396\,
            in1 => \N__29297\,
            in2 => \N__29285\,
            in3 => \N__48098\,
            lcout => n22019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i23_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35341\,
            in1 => \N__32002\,
            in2 => \N__29260\,
            in3 => \N__34425\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i24_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__34426\,
            in1 => \N__35343\,
            in2 => \N__29240\,
            in3 => \N__29256\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_303_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34960\,
            in2 => \_gnd_net_\,
            in3 => \N__35044\,
            lcout => n20590,
            ltout => \n20590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__30397\,
            in1 => \N__29238\,
            in2 => \N__30413\,
            in3 => \N__35344\,
            lcout => buf_adcdata_vac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_count_i0_i0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41437\,
            in2 => \N__30303\,
            in3 => \_gnd_net_\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => n19345,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30189\,
            in2 => \_gnd_net_\,
            in3 => \N__30170\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n19345,
            carryout => n19346,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30075\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n19346,
            carryout => n19347,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29973\,
            in2 => \_gnd_net_\,
            in3 => \N__29951\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n19347,
            carryout => n19348,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29859\,
            in2 => \_gnd_net_\,
            in3 => \N__29837\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n19348,
            carryout => n19349,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29757\,
            in2 => \_gnd_net_\,
            in3 => \N__29735\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n19349,
            carryout => n19350,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29649\,
            in2 => \_gnd_net_\,
            in3 => \N__29627\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n19350,
            carryout => n19351,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \N__29519\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n19351,
            carryout => n19352,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__41886\,
            sr => \N__41839\
        );

    \data_count_i0_i8_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30720\,
            in2 => \_gnd_net_\,
            in3 => \N__30698\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => n19353,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__41875\,
            sr => \N__41840\
        );

    \data_count_i0_i9_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30606\,
            in2 => \_gnd_net_\,
            in3 => \N__30695\,
            lcout => data_count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__41875\,
            sr => \N__41840\
        );

    \ADC_VAC.ADC_DATA_i8_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__30511\,
            in1 => \N__34624\,
            in2 => \N__35422\,
            in3 => \N__30584\,
            lcout => buf_adcdata_vac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_0_i19_3_lut_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56072\,
            in1 => \N__30545\,
            in2 => \_gnd_net_\,
            in3 => \N__30510\,
            lcout => n19_adj_1487,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i9_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34622\,
            in1 => \N__35394\,
            in2 => \N__30446\,
            in3 => \N__30823\,
            lcout => buf_adcdata_vac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i21_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30909\,
            in1 => \N__52990\,
            in2 => \N__51094\,
            in3 => \N__52076\,
            lcout => cmd_rdadctmp_21_adj_1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i10_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__30460\,
            in1 => \N__34623\,
            in2 => \N__30971\,
            in3 => \N__35395\,
            lcout => buf_adcdata_vac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_2_i19_3_lut_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56071\,
            in1 => \N__30497\,
            in2 => \_gnd_net_\,
            in3 => \N__30459\,
            lcout => n19_adj_1516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i18_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__30966\,
            in1 => \N__34430\,
            in2 => \N__30445\,
            in3 => \N__35396\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i19_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35393\,
            in1 => \N__30967\,
            in2 => \N__34518\,
            in3 => \N__34431\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i12_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__38148\,
            in1 => \N__51095\,
            in2 => \N__53156\,
            in3 => \N__52936\,
            lcout => buf_adcdata_iac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i13_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52933\,
            in1 => \N__53116\,
            in2 => \N__43578\,
            in3 => \N__30911\,
            lcout => buf_adcdata_iac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_5_i23_3_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30946\,
            in1 => \N__56236\,
            in2 => \_gnd_net_\,
            in3 => \N__38843\,
            lcout => n23_adj_1536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i22_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52935\,
            in1 => \N__30910\,
            in2 => \N__30876\,
            in3 => \N__52075\,
            lcout => cmd_rdadctmp_22_adj_1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54947\,
            in1 => \N__31009\,
            in2 => \N__49827\,
            in3 => \N__30895\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i14_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__52934\,
            in1 => \N__53117\,
            in2 => \N__30877\,
            in3 => \N__38352\,
            lcout => buf_adcdata_iac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i12_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49750\,
            in1 => \N__38972\,
            in2 => \N__44169\,
            in3 => \N__40326\,
            lcout => buf_dds0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_1_i19_3_lut_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56237\,
            in1 => \N__30854\,
            in2 => \_gnd_net_\,
            in3 => \N__30813\,
            lcout => n19_adj_1520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15012_3_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45916\,
            in1 => \N__31052\,
            in2 => \_gnd_net_\,
            in3 => \N__41728\,
            lcout => n17411,
            ltout => \n17411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15014_4_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__54888\,
            in1 => \N__49663\,
            in2 => \N__31169\,
            in3 => \N__31066\,
            lcout => \data_index_9_N_216_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__31067\,
            in1 => \N__31058\,
            in2 => \N__49758\,
            in3 => \N__54891\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__53586\,
            in1 => \N__48232\,
            in2 => \N__34864\,
            in3 => \N__49003\,
            lcout => n8828,
            ltout => \n8828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4419_3_lut_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41158\,
            in2 => \N__31034\,
            in3 => \N__31030\,
            lcout => n8_adj_1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i11_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__38555\,
            in1 => \N__40479\,
            in2 => \N__44309\,
            in3 => \N__38454\,
            lcout => buf_dds1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i13_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__30993\,
            in1 => \N__38556\,
            in2 => \N__47591\,
            in3 => \N__54890\,
            lcout => buf_dds1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__54889\,
            in1 => \N__39427\,
            in2 => \N__39449\,
            in3 => \N__49664\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_6_i16_3_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31275\,
            in1 => \N__31299\,
            in2 => \_gnd_net_\,
            in3 => \N__56244\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9341_1_lut_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50002\,
            lcout => n11757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i7_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__44586\,
            in1 => \N__38561\,
            in2 => \N__47681\,
            in3 => \N__38453\,
            lcout => buf_dds1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i6_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__31300\,
            in1 => \N__52507\,
            in2 => \N__49832\,
            in3 => \N__38954\,
            lcout => buf_dds0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i6_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__31276\,
            in1 => \N__38560\,
            in2 => \N__52511\,
            in3 => \N__38452\,
            lcout => buf_dds1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49767\,
            in1 => \N__49373\,
            in2 => \N__32371\,
            in3 => \N__43155\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57913\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_cnt_3774_3775__i1_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__31206\,
            in1 => \N__31245\,
            in2 => \_gnd_net_\,
            in3 => \N__31226\,
            lcout => wdtick_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32734\,
            ce => \N__31262\,
            sr => \N__40696\
        );

    \wdtick_cnt_3774_3775__i3_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010100000"
        )
    port map (
            in0 => \N__31228\,
            in1 => \_gnd_net_\,
            in2 => \N__31250\,
            in3 => \N__31207\,
            lcout => wdtick_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32734\,
            ce => \N__31262\,
            sr => \N__40696\
        );

    \wdtick_cnt_3774_3775__i2_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31244\,
            in2 => \_gnd_net_\,
            in3 => \N__31227\,
            lcout => wdtick_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32734\,
            ce => \N__31262\,
            sr => \N__40696\
        );

    \wdtick_flag_299_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__31249\,
            in1 => \N__31229\,
            in2 => \N__31211\,
            in3 => \N__49998\,
            lcout => wdtick_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32733\,
            ce => 'H',
            sr => \N__40697\
        );

    \SIG_DDS.tmp_buf_i0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__50178\,
            in1 => \N__50249\,
            in2 => \N__44728\,
            in3 => \N__31193\,
            lcout => \SIG_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57951\,
            ce => \N__31389\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19098_4_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100110"
        )
    port map (
            in0 => \N__50248\,
            in1 => \N__50366\,
            in2 => \N__44811\,
            in3 => \N__50177\,
            lcout => \SIG_DDS.n12738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15029_2_lut_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35716\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31369\,
            lcout => \OUT_SYNCCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0off_i0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32609\,
            in2 => \_gnd_net_\,
            in3 => \N__31334\,
            lcout => \ADC_VDC.genclk.t0off_0\,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \ADC_VDC.genclk.n19468\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i1_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32579\,
            in2 => \N__57324\,
            in3 => \N__31331\,
            lcout => \ADC_VDC.genclk.t0off_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19468\,
            carryout => \ADC_VDC.genclk.n19469\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i2_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57251\,
            in2 => \N__31328\,
            in3 => \N__31313\,
            lcout => \ADC_VDC.genclk.t0off_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19469\,
            carryout => \ADC_VDC.genclk.n19470\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i3_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32678\,
            in2 => \N__57325\,
            in3 => \N__31310\,
            lcout => \ADC_VDC.genclk.t0off_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19470\,
            carryout => \ADC_VDC.genclk.n19471\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i4_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57255\,
            in2 => \N__32597\,
            in3 => \N__31307\,
            lcout => \ADC_VDC.genclk.t0off_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19471\,
            carryout => \ADC_VDC.genclk.n19472\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i5_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32665\,
            in2 => \N__57326\,
            in3 => \N__31304\,
            lcout => \ADC_VDC.genclk.t0off_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19472\,
            carryout => \ADC_VDC.genclk.n19473\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i6_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57259\,
            in2 => \N__32624\,
            in3 => \N__31475\,
            lcout => \ADC_VDC.genclk.t0off_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19473\,
            carryout => \ADC_VDC.genclk.n19474\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i7_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31471\,
            in2 => \N__57327\,
            in3 => \N__31457\,
            lcout => \ADC_VDC.genclk.t0off_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19474\,
            carryout => \ADC_VDC.genclk.n19475\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__31601\,
            sr => \N__33880\
        );

    \ADC_VDC.genclk.t0off_i8_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32651\,
            in2 => \N__57384\,
            in3 => \N__31454\,
            lcout => \ADC_VDC.genclk.t0off_8\,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => \ADC_VDC.genclk.n19476\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i9_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57346\,
            in2 => \N__32549\,
            in3 => \N__31451\,
            lcout => \ADC_VDC.genclk.t0off_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19476\,
            carryout => \ADC_VDC.genclk.n19477\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i10_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31448\,
            in2 => \N__57381\,
            in3 => \N__31436\,
            lcout => \ADC_VDC.genclk.t0off_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19477\,
            carryout => \ADC_VDC.genclk.n19478\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i11_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57334\,
            in2 => \N__32519\,
            in3 => \N__31433\,
            lcout => \ADC_VDC.genclk.t0off_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19478\,
            carryout => \ADC_VDC.genclk.n19479\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i12_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31430\,
            in2 => \N__57382\,
            in3 => \N__31418\,
            lcout => \ADC_VDC.genclk.t0off_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19479\,
            carryout => \ADC_VDC.genclk.n19480\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i13_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57338\,
            in2 => \N__32693\,
            in3 => \N__31415\,
            lcout => \ADC_VDC.genclk.t0off_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19480\,
            carryout => \ADC_VDC.genclk.n19481\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i14_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32561\,
            in2 => \N__57383\,
            in3 => \N__31412\,
            lcout => \ADC_VDC.genclk.t0off_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19481\,
            carryout => \ADC_VDC.genclk.n19482\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \ADC_VDC.genclk.t0off_i15_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32533\,
            in1 => \N__57342\,
            in2 => \_gnd_net_\,
            in3 => \N__31604\,
            lcout => \ADC_VDC.genclk.t0off_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__31597\,
            sr => \N__33872\
        );

    \i19_4_lut_adj_249_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100010001"
        )
    port map (
            in0 => \N__54174\,
            in1 => \N__37516\,
            in2 => \N__54383\,
            in3 => \N__31625\,
            lcout => OPEN,
            ltout => \n12_adj_1615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_250_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42785\,
            in2 => \N__31577\,
            in3 => \N__50926\,
            lcout => n12236,
            ltout => \n12236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12388_2_lut_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31574\,
            in3 => \N__54911\,
            lcout => n14801,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50776\,
            in1 => \N__31571\,
            in2 => \_gnd_net_\,
            in3 => \N__54177\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57806\,
            ce => \N__31489\,
            sr => \N__31669\
        );

    \comm_buf_5__i1_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54175\,
            in1 => \N__45365\,
            in2 => \_gnd_net_\,
            in3 => \N__31556\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57806\,
            ce => \N__31489\,
            sr => \N__31669\
        );

    \comm_buf_5__i2_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47241\,
            in1 => \N__31538\,
            in2 => \_gnd_net_\,
            in3 => \N__54178\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57806\,
            ce => \N__31489\,
            sr => \N__31669\
        );

    \comm_buf_5__i3_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54176\,
            in1 => \N__40776\,
            in2 => \_gnd_net_\,
            in3 => \N__31523\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57806\,
            ce => \N__31489\,
            sr => \N__31669\
        );

    \comm_buf_5__i4_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40645\,
            in1 => \N__31508\,
            in2 => \_gnd_net_\,
            in3 => \N__54179\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57806\,
            ce => \N__31489\,
            sr => \N__31669\
        );

    \mux_143_Mux_4_i2_3_lut_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36986\,
            in1 => \N__31823\,
            in2 => \_gnd_net_\,
            in3 => \N__54382\,
            lcout => OPEN,
            ltout => \n2_adj_1587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__50687\,
            in1 => \N__31631\,
            in2 => \N__31655\,
            in3 => \N__31637\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57808\,
            ce => \N__46223\,
            sr => \N__46140\
        );

    \i18721_2_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31904\,
            in2 => \_gnd_net_\,
            in3 => \N__54379\,
            lcout => n21324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_4_i4_3_lut_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54380\,
            in1 => \N__31652\,
            in2 => \_gnd_net_\,
            in3 => \N__37721\,
            lcout => OPEN,
            ltout => \n4_adj_1588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19504_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__31646\,
            in1 => \N__50554\,
            in2 => \N__31640\,
            in3 => \N__50686\,
            lcout => n22136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_4_i1_3_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54381\,
            in1 => \N__51182\,
            in2 => \_gnd_net_\,
            in3 => \N__44120\,
            lcout => n1_adj_1586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50553\,
            in2 => \N__43070\,
            in3 => \N__50685\,
            lcout => n19006,
            ltout => \n19006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_246_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__54378\,
            in1 => \N__54150\,
            in2 => \N__31619\,
            in3 => \N__37517\,
            lcout => n12_adj_1639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i7_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54166\,
            in1 => \N__51393\,
            in2 => \_gnd_net_\,
            in3 => \N__31616\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \comm_buf_2__i6_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40234\,
            in1 => \N__31862\,
            in2 => \_gnd_net_\,
            in3 => \N__54168\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \comm_buf_2__i5_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54165\,
            in1 => \N__51043\,
            in2 => \_gnd_net_\,
            in3 => \N__31850\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \comm_buf_2__i4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54139\,
            in1 => \N__31838\,
            in2 => \_gnd_net_\,
            in3 => \N__40646\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \comm_buf_2__i3_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54164\,
            in1 => \N__40793\,
            in2 => \_gnd_net_\,
            in3 => \N__31817\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \comm_buf_2__i2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47242\,
            in1 => \N__31805\,
            in2 => \_gnd_net_\,
            in3 => \N__54167\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57813\,
            ce => \N__34217\,
            sr => \N__34190\
        );

    \ADC_VDC.cmd_rdadctmp_i23_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__31793\,
            in1 => \N__31763\,
            in2 => \N__31744\,
            in3 => \N__32869\,
            lcout => \ADC_VDC.cmd_rdadctmp_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40131\,
            ce => \N__31724\,
            sr => \N__31718\
        );

    \RTD.i2_3_lut_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33766\,
            in1 => \N__33789\,
            in2 => \_gnd_net_\,
            in3 => \N__33806\,
            lcout => \RTD.n17720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_6_i23_3_lut_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45017\,
            in1 => \N__56106\,
            in2 => \_gnd_net_\,
            in3 => \N__32372\,
            lcout => n23_adj_1534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__32100\,
            in1 => \N__32027\,
            in2 => \N__40569\,
            in3 => \N__51405\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22160_bdd_4_lut_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000100010"
        )
    port map (
            in0 => \N__31966\,
            in1 => \N__48094\,
            in2 => \N__31928\,
            in3 => \N__31913\,
            lcout => n22163,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i20_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__34519\,
            in1 => \N__34410\,
            in2 => \N__34686\,
            in3 => \N__35376\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__37618\,
            in1 => \N__54907\,
            in2 => \N__40801\,
            in3 => \N__51312\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i4_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__51313\,
            in1 => \N__31903\,
            in2 => \N__54962\,
            in3 => \N__40654\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18755_2_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53561\,
            in2 => \_gnd_net_\,
            in3 => \N__31889\,
            lcout => n20962,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__48816\,
            in1 => \N__32121\,
            in2 => \N__47252\,
            in3 => \N__32032\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__47998\,
            in1 => \N__45377\,
            in2 => \N__32044\,
            in3 => \N__32120\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i22_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35406\,
            in1 => \N__34702\,
            in2 => \N__32003\,
            in3 => \N__34428\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__47997\,
            in1 => \N__55816\,
            in2 => \_gnd_net_\,
            in3 => \N__48815\,
            lcout => n10733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i21_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35405\,
            in1 => \N__34701\,
            in2 => \N__34687\,
            in3 => \N__34427\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i17_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34594\,
            in1 => \N__35408\,
            in2 => \N__34487\,
            in3 => \N__43947\,
            lcout => buf_adcdata_vac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__55817\,
            in1 => \N__50783\,
            in2 => \N__32123\,
            in3 => \N__32028\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i14_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__35407\,
            in2 => \N__38077\,
            in3 => \N__32001\,
            lcout => buf_adcdata_vac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__46547\,
            in1 => \N__54803\,
            in2 => \N__41234\,
            in3 => \N__31985\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => n19393,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__46816\,
            in1 => \N__54807\,
            in2 => \N__43421\,
            in3 => \N__31982\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n19393,
            carryout => n19394,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__44054\,
            in1 => \N__54804\,
            in2 => \N__46870\,
            in3 => \N__31979\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n19394,
            carryout => n19395,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47843\,
            in1 => \N__54808\,
            in2 => \N__37880\,
            in3 => \N__31976\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n19395,
            carryout => n19396,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__51119\,
            in1 => \N__54805\,
            in2 => \N__38218\,
            in3 => \N__31973\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n19396,
            carryout => n19397,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47322\,
            in1 => \N__54809\,
            in2 => \N__43489\,
            in3 => \N__31970\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n19397,
            carryout => n19398,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__52175\,
            in1 => \N__54806\,
            in2 => \N__37786\,
            in3 => \N__32174\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n19398,
            carryout => n19399,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47606\,
            in1 => \N__54810\,
            in2 => \N__49249\,
            in3 => \N__32171\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n19399,
            carryout => n19400,
            clk => \N__57839\,
            ce => \N__39061\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__44478\,
            in1 => \N__54892\,
            in2 => \N__41584\,
            in3 => \N__32168\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => n19401,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47462\,
            in1 => \N__54899\,
            in2 => \N__44347\,
            in3 => \N__32165\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n19401,
            carryout => n19402,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__39313\,
            in1 => \N__54893\,
            in2 => \N__34165\,
            in3 => \N__32162\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n19402,
            carryout => n19403,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__39274\,
            in1 => \N__54900\,
            in2 => \N__40864\,
            in3 => \N__32159\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n19403,
            carryout => n19404,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__44077\,
            in1 => \N__54894\,
            in2 => \N__40945\,
            in3 => \N__32156\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n19404,
            carryout => n19405,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__47587\,
            in1 => \N__54901\,
            in2 => \N__32149\,
            in3 => \N__32129\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n19405,
            carryout => n19406,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__39190\,
            in1 => \N__54895\,
            in2 => \N__36274\,
            in3 => \N__32126\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n19406,
            carryout => n19407,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46795\,
            in1 => \N__32267\,
            in2 => \N__54960\,
            in3 => \N__32291\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57849\,
            ce => \N__39065\,
            sr => \_gnd_net_\
        );

    \i18129_4_lut_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__36715\,
            in1 => \N__36418\,
            in2 => \N__41050\,
            in3 => \N__36335\,
            lcout => n20742,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22166_bdd_4_lut_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__49011\,
            in1 => \N__41303\,
            in2 => \N__47765\,
            in3 => \N__32240\,
            lcout => OPEN,
            ltout => \n22169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1545458_i1_3_lut_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__48714\,
            in1 => \_gnd_net_\,
            in2 => \N__32288\,
            in3 => \N__32285\,
            lcout => n30_adj_1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19099_4_lut_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100110011"
        )
    port map (
            in0 => \N__36419\,
            in1 => \N__36716\,
            in2 => \N__36062\,
            in3 => \N__41035\,
            lcout => OPEN,
            ltout => \n20568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_309_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__36717\,
            in1 => \N__32255\,
            in2 => \N__32270\,
            in3 => \N__36336\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_end_309C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i26_3_lut_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32266\,
            in1 => \N__56073\,
            in2 => \_gnd_net_\,
            in3 => \N__32254\,
            lcout => OPEN,
            ltout => \n26_adj_1528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19523_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__55586\,
            in1 => \N__48228\,
            in2 => \N__32243\,
            in3 => \N__49010\,
            lcout => n22166,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_310_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__41036\,
            in1 => \N__36718\,
            in2 => \N__32217\,
            in3 => \N__32234\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_end_309C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14176_4_lut_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__41626\,
            in1 => \N__43925\,
            in2 => \N__36725\,
            in3 => \N__36191\,
            lcout => OPEN,
            ltout => \n16594_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000010001"
        )
    port map (
            in0 => \N__36416\,
            in1 => \N__36724\,
            in2 => \N__32309\,
            in3 => \N__32306\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__36146\,
            sr => \N__36352\
        );

    \eis_state_1__bdd_4_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__35885\,
            in1 => \N__36415\,
            in2 => \N__35897\,
            in3 => \N__41021\,
            lcout => n22196,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_197_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__41625\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36190\,
            lcout => n16602,
            ltout => \n16602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__36417\,
            in1 => \N__41023\,
            in2 => \N__32300\,
            in3 => \N__35432\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__36146\,
            sr => \N__36352\
        );

    \i34_3_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36414\,
            in1 => \N__41433\,
            in2 => \_gnd_net_\,
            in3 => \N__32297\,
            lcout => n13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_168_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__32483\,
            in2 => \N__38995\,
            in3 => \N__32337\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__41284\,
            in1 => \N__49691\,
            in2 => \N__41167\,
            in3 => \N__49371\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__49368\,
            in1 => \N__44155\,
            in2 => \N__49775\,
            in3 => \N__38994\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32426\,
            in1 => \N__32465\,
            in2 => \N__42438\,
            in3 => \N__32361\,
            lcout => n23_adj_1624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__49367\,
            in1 => \N__42987\,
            in2 => \N__49774\,
            in3 => \N__32338\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__44308\,
            in1 => \N__49369\,
            in2 => \N__42439\,
            in3 => \N__49698\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_176_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__38014\,
            in1 => \N__32320\,
            in2 => \N__32393\,
            in3 => \N__41283\,
            lcout => n17_adj_1612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__45911\,
            in1 => \N__49370\,
            in2 => \N__43528\,
            in3 => \N__49699\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41432\,
            in2 => \N__32324\,
            in3 => \_gnd_net_\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => n19369,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__36627\,
            sr => \N__36446\
        );

    \add_79_2_THRU_CRY_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57410\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n19369,
            carryout => \n19369_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__57423\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_0_THRU_CO\,
            carryout => \n19369_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_2_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57414\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_1_THRU_CO\,
            carryout => \n19369_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_3_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__57424\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_2_THRU_CO\,
            carryout => \n19369_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_4_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57418\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_3_THRU_CO\,
            carryout => \n19369_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_5_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__57425\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_4_THRU_CO\,
            carryout => \n19369_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_79_2_THRU_CRY_6_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57422\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19369_THRU_CRY_5_THRU_CO\,
            carryout => \n19369_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38809\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => n19370,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39235\,
            in2 => \_gnd_net_\,
            in3 => \N__32405\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n19370,
            carryout => n19371,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36235\,
            in2 => \_gnd_net_\,
            in3 => \N__32402\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n19371,
            carryout => n19372,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38788\,
            in2 => \_gnd_net_\,
            in3 => \N__32399\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n19372,
            carryout => n19373,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i5_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36253\,
            in2 => \_gnd_net_\,
            in3 => \N__32396\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n19373,
            carryout => n19374,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i6_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32389\,
            in2 => \_gnd_net_\,
            in3 => \N__32375\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n19374,
            carryout => n19375,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i7_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39253\,
            in2 => \_gnd_net_\,
            in3 => \N__32492\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n19375,
            carryout => n19376,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i8_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36217\,
            in2 => \_gnd_net_\,
            in3 => \N__32489\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n19376,
            carryout => n19377,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__36635\,
            sr => \N__36598\
        );

    \acadc_skipcnt_i0_i9_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36481\,
            in2 => \_gnd_net_\,
            in3 => \N__32486\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => n19378,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i10_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32482\,
            in2 => \_gnd_net_\,
            in3 => \N__32468\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n19378,
            carryout => n19379,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i11_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32464\,
            in2 => \_gnd_net_\,
            in3 => \N__32450\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n19379,
            carryout => n19380,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i12_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32446\,
            in2 => \_gnd_net_\,
            in3 => \N__32432\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n19380,
            carryout => n19381,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i13_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38857\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n19381,
            carryout => n19382,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i14_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32425\,
            in2 => \_gnd_net_\,
            in3 => \N__32411\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n19382,
            carryout => n19383,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \acadc_skipcnt_i0_i15_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36496\,
            in2 => \_gnd_net_\,
            in3 => \N__32744\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__36634\,
            sr => \N__36599\
        );

    \SecClk_302_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39746\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__32677\,
            in2 => \N__32666\,
            in3 => \N__32650\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i18779_4_lut_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32504\,
            in1 => \N__32639\,
            in2 => \N__32630\,
            in3 => \N__32567\,
            lcout => \ADC_VDC.genclk.n21206\,
            ltout => \ADC_VDC.genclk.n21206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i0_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__33673\,
            in1 => \N__40170\,
            in2 => \N__32627\,
            in3 => \N__37216\,
            lcout => \ADC_VDC.genclk.div_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19076_4_lut_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__32620\,
            in1 => \N__32608\,
            in2 => \N__32596\,
            in3 => \N__32578\,
            lcout => \ADC_VDC.genclk.n21208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32560\,
            in1 => \N__32545\,
            in2 => \N__32534\,
            in3 => \N__32515\,
            lcout => \ADC_VDC.genclk.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19182_2_lut_4_lut_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011111111111"
        )
    port map (
            in0 => \N__40162\,
            in1 => \N__32498\,
            in2 => \N__37217\,
            in3 => \N__33668\,
            lcout => \ADC_VDC.genclk.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i1_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33669\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40163\,
            lcout => \ADC_VDC.genclk.div_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i1C_net\,
            ce => \N__33686\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12662_2_lut_2_lut_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__40160\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33667\,
            lcout => \ADC_VDC.genclk.n15067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.genclk.div_state_1__N_1275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16075_4_lut_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010111010"
        )
    port map (
            in0 => \N__33300\,
            in1 => \N__33097\,
            in2 => \N__33383\,
            in3 => \N__32895\,
            lcout => \ADC_VDC.n11766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_39_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__33630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33524\,
            lcout => \ADC_VDC.n62\,
            ltout => \ADC_VDC.n62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i24_4_lut_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010111010"
        )
    port map (
            in0 => \N__33299\,
            in1 => \N__33096\,
            in2 => \N__32909\,
            in3 => \N__32894\,
            lcout => \ADC_VDC.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0on_i0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37232\,
            in2 => \_gnd_net_\,
            in3 => \N__32753\,
            lcout => \ADC_VDC.genclk.t0on_0\,
            ltout => OPEN,
            carryin => \bfn_13_5_0_\,
            carryout => \ADC_VDC.genclk.n19483\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i1_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37265\,
            in2 => \N__57388\,
            in3 => \N__32750\,
            lcout => \ADC_VDC.genclk.t0on_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19483\,
            carryout => \ADC_VDC.genclk.n19484\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i2_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57353\,
            in2 => \N__37064\,
            in3 => \N__32747\,
            lcout => \ADC_VDC.genclk.t0on_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19484\,
            carryout => \ADC_VDC.genclk.n19485\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i3_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37187\,
            in2 => \N__57389\,
            in3 => \N__33713\,
            lcout => \ADC_VDC.genclk.t0on_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19485\,
            carryout => \ADC_VDC.genclk.n19486\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i4_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57357\,
            in2 => \N__37252\,
            in3 => \N__33710\,
            lcout => \ADC_VDC.genclk.t0on_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19486\,
            carryout => \ADC_VDC.genclk.n19487\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i5_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37174\,
            in2 => \N__57390\,
            in3 => \N__33707\,
            lcout => \ADC_VDC.genclk.t0on_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19487\,
            carryout => \ADC_VDC.genclk.n19488\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i6_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57361\,
            in2 => \N__37280\,
            in3 => \N__33704\,
            lcout => \ADC_VDC.genclk.t0on_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19488\,
            carryout => \ADC_VDC.genclk.n19489\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i7_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37048\,
            in2 => \N__57391\,
            in3 => \N__33701\,
            lcout => \ADC_VDC.genclk.t0on_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19489\,
            carryout => \ADC_VDC.genclk.n19490\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__33908\,
            sr => \N__33881\
        );

    \ADC_VDC.genclk.t0on_i8_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57375\,
            in2 => \N__37160\,
            in3 => \N__33698\,
            lcout => \ADC_VDC.genclk.t0on_8\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \ADC_VDC.genclk.n19491\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i9_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37124\,
            in2 => \N__57394\,
            in3 => \N__33695\,
            lcout => \ADC_VDC.genclk.t0on_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19491\,
            carryout => \ADC_VDC.genclk.n19492\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i10_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57365\,
            in2 => \N__37034\,
            in3 => \N__33692\,
            lcout => \ADC_VDC.genclk.t0on_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19492\,
            carryout => \ADC_VDC.genclk.n19493\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i11_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37097\,
            in2 => \N__57392\,
            in3 => \N__33689\,
            lcout => \ADC_VDC.genclk.t0on_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19493\,
            carryout => \ADC_VDC.genclk.n19494\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i12_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57369\,
            in2 => \N__37079\,
            in3 => \N__33920\,
            lcout => \ADC_VDC.genclk.t0on_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19494\,
            carryout => \ADC_VDC.genclk.n19495\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i13_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37199\,
            in2 => \N__57393\,
            in3 => \N__33917\,
            lcout => \ADC_VDC.genclk.t0on_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19495\,
            carryout => \ADC_VDC.genclk.n19496\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i14_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57373\,
            in2 => \N__37139\,
            in3 => \N__33914\,
            lcout => \ADC_VDC.genclk.t0on_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19496\,
            carryout => \ADC_VDC.genclk.n19497\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \ADC_VDC.genclk.t0on_i15_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57374\,
            in1 => \N__37111\,
            in2 => \_gnd_net_\,
            in3 => \N__33911\,
            lcout => \ADC_VDC.genclk.t0on_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__33907\,
            sr => \N__33873\
        );

    \RTD.bit_cnt_3782__i3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__33809\,
            in1 => \N__33823\,
            in2 => \N__33776\,
            in3 => \N__33791\,
            lcout => \RTD.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43735\,
            ce => \N__33749\,
            sr => \N__33731\
        );

    \RTD.bit_cnt_3782__i1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33768\,
            in2 => \_gnd_net_\,
            in3 => \N__33807\,
            lcout => \RTD.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43735\,
            ce => \N__33749\,
            sr => \N__33731\
        );

    \RTD.bit_cnt_3782__i2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__33808\,
            in1 => \_gnd_net_\,
            in2 => \N__33775\,
            in3 => \N__33790\,
            lcout => \RTD.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43735\,
            ce => \N__33749\,
            sr => \N__33731\
        );

    \RTD.bit_cnt_3782__i0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33767\,
            lcout => \RTD.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__43735\,
            ce => \N__33749\,
            sr => \N__33731\
        );

    \i1_3_lut_adj_245_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__42783\,
            in1 => \N__50931\,
            in2 => \_gnd_net_\,
            in3 => \N__37478\,
            lcout => n12152,
            ltout => \n12152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12374_2_lut_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34085\,
            in3 => \N__54829\,
            lcout => n14787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_247_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__42784\,
            in1 => \_gnd_net_\,
            in2 => \N__34082\,
            in3 => \N__50930\,
            lcout => n12194,
            ltout => \n12194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12381_2_lut_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34073\,
            in3 => \N__54828\,
            lcout => n14794,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_0_i22_3_lut_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34063\,
            in1 => \N__33926\,
            in2 => \_gnd_net_\,
            in3 => \N__49074\,
            lcout => OPEN,
            ltout => \n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_136_Mux_0_i30_3_lut_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48738\,
            in1 => \_gnd_net_\,
            in2 => \N__34037\,
            in3 => \N__34034\,
            lcout => OPEN,
            ltout => \n30_adj_1484_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i0_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50778\,
            in2 => \N__34022\,
            in3 => \N__53842\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57823\,
            ce => \N__34216\,
            sr => \N__34189\
        );

    \mux_136_Mux_1_i30_3_lut_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48739\,
            in1 => \_gnd_net_\,
            in2 => \N__34019\,
            in3 => \N__34004\,
            lcout => OPEN,
            ltout => \n30_adj_1504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i1_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__45364\,
            in1 => \_gnd_net_\,
            in2 => \N__33989\,
            in3 => \N__53843\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57823\,
            ce => \N__34216\,
            sr => \N__34189\
        );

    \mux_136_Mux_0_i19_3_lut_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33986\,
            in1 => \N__33965\,
            in2 => \_gnd_net_\,
            in3 => \N__56143\,
            lcout => n19_adj_1485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_242_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__53566\,
            in1 => \N__42782\,
            in2 => \N__50933\,
            in3 => \N__37793\,
            lcout => n12110,
            ltout => \n12110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12367_2_lut_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34193\,
            in3 => \N__54735\,
            lcout => n14780,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18291_3_lut_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55948\,
            in1 => \N__34166\,
            in2 => \_gnd_net_\,
            in3 => \N__42068\,
            lcout => OPEN,
            ltout => \n20905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19514_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__48217\,
            in1 => \N__34091\,
            in2 => \N__34145\,
            in3 => \N__48875\,
            lcout => OPEN,
            ltout => \n22148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22148_bdd_4_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48876\,
            in1 => \N__34142\,
            in2 => \N__34127\,
            in3 => \N__34715\,
            lcout => OPEN,
            ltout => \n22151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18275_3_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34124\,
            in2 => \N__34112\,
            in3 => \N__48619\,
            lcout => OPEN,
            ltout => \n20889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i2_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47247\,
            in2 => \N__34109\,
            in3 => \N__54089\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57832\,
            ce => \N__42725\,
            sr => \N__42856\
        );

    \i18735_2_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34106\,
            in2 => \_gnd_net_\,
            in3 => \N__55947\,
            lcout => n20906,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_i8_2_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__48874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48216\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_278_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__48215\,
            in1 => \N__55946\,
            in2 => \N__34838\,
            in3 => \N__48873\,
            lcout => n20672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i1_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34650\,
            in1 => \N__35404\,
            in2 => \N__34772\,
            in3 => \N__34734\,
            lcout => buf_adcdata_vac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18226_3_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55945\,
            in1 => \N__35678\,
            in2 => \_gnd_net_\,
            in3 => \N__42017\,
            lcout => n20840,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i13_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34649\,
            in1 => \N__35403\,
            in2 => \N__34706\,
            in3 => \N__46635\,
            lcout => buf_adcdata_vac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i12_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__35400\,
            in1 => \N__34651\,
            in2 => \N__34688\,
            in3 => \N__35593\,
            lcout => buf_adcdata_vac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i11_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34648\,
            in1 => \N__35402\,
            in2 => \N__38290\,
            in3 => \N__34520\,
            lcout => buf_adcdata_vac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i26_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35401\,
            in1 => \N__34483\,
            in2 => \N__34234\,
            in3 => \N__34429\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i39_3_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__48090\,
            in1 => \N__55944\,
            in2 => \_gnd_net_\,
            in3 => \N__48856\,
            lcout => OPEN,
            ltout => \n24_adj_1622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i41_3_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48703\,
            in2 => \N__35630\,
            in3 => \N__36572\,
            lcout => n21_adj_1618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_4_i19_3_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35627\,
            in1 => \N__35589\,
            in2 => \_gnd_net_\,
            in3 => \N__55949\,
            lcout => n19_adj_1509,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_214_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41051\,
            in2 => \_gnd_net_\,
            in3 => \N__36432\,
            lcout => OPEN,
            ltout => \n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3798_3_lut_3_lut_4_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__41418\,
            in1 => \N__36719\,
            in2 => \N__35573\,
            in3 => \N__36337\,
            lcout => \iac_raw_buf_N_735\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101001011000"
        )
    port map (
            in0 => \N__36720\,
            in1 => \N__41052\,
            in2 => \N__36437\,
            in3 => \N__41419\,
            lcout => n17_adj_1645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.DTRIG_39_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__35416\,
            in1 => \N__35048\,
            in2 => \N__34967\,
            in3 => \N__36118\,
            lcout => acadc_dtrig_v,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_340_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41623\,
            in1 => \N__43878\,
            in2 => \_gnd_net_\,
            in3 => \N__41493\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__54823\,
            in1 => \N__53567\,
            in2 => \N__34877\,
            in3 => \N__34865\,
            lcout => n10534,
            ltout => \n10534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \auxmode_337_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44281\,
            in1 => \_gnd_net_\,
            in2 => \N__34841\,
            in3 => \N__35698\,
            lcout => auxmode,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14180_1_lut_2_lut_3_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__36085\,
            in1 => \_gnd_net_\,
            in2 => \N__36122\,
            in3 => \N__36675\,
            lcout => n16598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36111\,
            in2 => \_gnd_net_\,
            in3 => \N__36083\,
            lcout => \iac_raw_buf_N_737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18743_2_lut_3_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__36084\,
            in1 => \_gnd_net_\,
            in2 => \N__36121\,
            in3 => \N__36676\,
            lcout => n20957,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.DTRIG_39_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__35876\,
            in1 => \N__35804\,
            in2 => \N__53001\,
            in3 => \N__36086\,
            lcout => acadc_dtrig_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ICE_GPMO_0_I_0_3_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35741\,
            in1 => \N__35697\,
            in2 => \_gnd_net_\,
            in3 => \N__35673\,
            lcout => acadc_rst,
            ltout => \acadc_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_4_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__36674\,
            in1 => \N__41045\,
            in2 => \N__35681\,
            in3 => \N__36421\,
            lcout => n13473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tacadc_rst_338_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42970\,
            in1 => \N__43879\,
            in2 => \_gnd_net_\,
            in3 => \N__35674\,
            lcout => tacadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18184_3_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35660\,
            in1 => \N__35642\,
            in2 => \_gnd_net_\,
            in3 => \N__48335\,
            lcout => n20798,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_201_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__41624\,
            in1 => \N__36128\,
            in2 => \N__36431\,
            in3 => \N__44905\,
            lcout => OPEN,
            ltout => \n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19147_3_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41020\,
            in2 => \N__36158\,
            in3 => \N__36685\,
            lcout => n11760,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18865_2_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__43920\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36420\,
            lcout => OPEN,
            ltout => \n21099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__41022\,
            in1 => \N__36686\,
            in2 => \N__36155\,
            in3 => \N__36152\,
            lcout => \eis_end_N_725\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i2C_net\,
            ce => \N__36142\,
            sr => \N__36338\
        );

    \i15032_2_lut_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36119\,
            in2 => \_gnd_net_\,
            in3 => \N__36081\,
            lcout => n17430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_263_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36120\,
            in2 => \N__43924\,
            in3 => \N__36082\,
            lcout => n4_adj_1569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36023\,
            in1 => \N__54967\,
            in2 => \N__49780\,
            in3 => \N__36014\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6444_3_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41747\,
            in1 => \N__37970\,
            in2 => \_gnd_net_\,
            in3 => \N__36039\,
            lcout => n8_adj_1563,
            ltout => \n8_adj_1563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_3_i15_4_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49708\,
            in1 => \N__54966\,
            in2 => \N__36017\,
            in3 => \N__36013\,
            lcout => \data_index_9_N_216_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__49343\,
            in1 => \N__49709\,
            in2 => \N__37930\,
            in3 => \N__37971\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49710\,
            in1 => \N__49342\,
            in2 => \N__41656\,
            in3 => \N__41494\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36254\,
            in1 => \N__36239\,
            in2 => \N__37929\,
            in3 => \N__43524\,
            lcout => OPEN,
            ltout => \n20_adj_1617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__36221\,
            in1 => \N__41646\,
            in2 => \N__36203\,
            in3 => \N__38819\,
            lcout => OPEN,
            ltout => \n26_adj_1640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_179_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38774\,
            in1 => \N__36200\,
            in2 => \N__36194\,
            in3 => \N__36452\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6434_3_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51168\,
            in1 => \N__38755\,
            in2 => \_gnd_net_\,
            in3 => \N__41729\,
            lcout => n8_adj_1561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__49357\,
            in1 => \N__49686\,
            in2 => \N__52506\,
            in3 => \N__38013\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__44608\,
            in1 => \N__45556\,
            in2 => \N__49773\,
            in3 => \N__49359\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__49358\,
            in1 => \N__49687\,
            in2 => \N__47673\,
            in3 => \N__49176\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6454_3_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36180\,
            in1 => \N__47139\,
            in2 => \_gnd_net_\,
            in3 => \N__41730\,
            lcout => n8_adj_1565,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__36500\,
            in1 => \N__36482\,
            in2 => \N__47787\,
            in3 => \N__44607\,
            lcout => OPEN,
            ltout => \n24_adj_1537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39221\,
            in1 => \N__36467\,
            in2 => \N__36461\,
            in3 => \N__36458\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19175_2_lut_3_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36345\,
            in1 => \N__41049\,
            in2 => \_gnd_net_\,
            in3 => \N__36708\,
            lcout => n20789,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i5_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__36295\,
            in1 => \N__38567\,
            in2 => \N__47327\,
            in3 => \N__54847\,
            lcout => buf_dds1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i7_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__38950\,
            in1 => \N__49720\,
            in2 => \N__47680\,
            in3 => \N__44562\,
            lcout => buf_dds0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19179_3_lut_4_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__36707\,
            in1 => \N__36433\,
            in2 => \N__41054\,
            in3 => \N__36344\,
            lcout => n11670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_5_i16_3_lut_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36291\,
            in1 => \N__36547\,
            in2 => \_gnd_net_\,
            in3 => \N__56298\,
            lcout => n16_adj_1496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12224_12225_set_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55400\,
            in1 => \N__55373\,
            in2 => \_gnd_net_\,
            in3 => \N__55349\,
            lcout => \comm_spi.n14642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57035\,
            ce => 'H',
            sr => \N__41930\
        );

    \i19065_2_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36275\,
            in2 => \_gnd_net_\,
            in3 => \N__56340\,
            lcout => n21037,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19118_2_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36709\,
            in2 => \_gnd_net_\,
            in3 => \N__36617\,
            lcout => n14687,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_237_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36586\,
            in2 => \_gnd_net_\,
            in3 => \N__46581\,
            lcout => n10713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39886\,
            in1 => \N__39709\,
            in2 => \N__39575\,
            in3 => \N__39511\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i5_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49781\,
            in1 => \N__36543\,
            in2 => \N__45917\,
            in3 => \N__38966\,
            lcout => buf_dds0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18827_2_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__42041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56363\,
            lcout => n21067,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_174_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39496\,
            in1 => \N__39610\,
            in2 => \N__39680\,
            in3 => \N__39541\,
            lcout => OPEN,
            ltout => \n27_adj_1551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36977\,
            in1 => \N__36506\,
            in2 => \N__36524\,
            in3 => \N__36521\,
            lcout => OPEN,
            ltout => \n19608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_187_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__39808\,
            in1 => \N__36971\,
            in2 => \N__36515\,
            in3 => \N__36512\,
            lcout => n14731,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_175_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => n10_adj_1594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_173_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39871\,
            in1 => \N__39724\,
            in2 => \N__39629\,
            in3 => \N__39556\,
            lcout => n26_adj_1543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_172_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39526\,
            in1 => \N__39589\,
            in2 => \N__39842\,
            in3 => \N__39661\,
            lcout => n28_adj_1621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_177_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39793\,
            in1 => \N__39823\,
            in2 => \N__39647\,
            in3 => \N__39775\,
            lcout => n14_adj_1592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22112_bdd_4_lut_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48362\,
            in1 => \N__36965\,
            in2 => \N__36926\,
            in3 => \N__36779\,
            lcout => OPEN,
            ltout => \n22115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18242_3_lut_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49118\,
            in2 => \N__36887\,
            in3 => \N__36884\,
            lcout => n20856,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19509_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__36865\,
            in1 => \N__48361\,
            in2 => \N__36824\,
            in3 => \N__56299\,
            lcout => n22112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19439_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__48363\,
            in1 => \N__42629\,
            in2 => \N__36773\,
            in3 => \N__49119\,
            lcout => OPEN,
            ltout => \n22070_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22070_bdd_4_lut_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49120\,
            in1 => \N__36752\,
            in2 => \N__36737\,
            in3 => \N__39170\,
            lcout => OPEN,
            ltout => \n22073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1544855_i1_3_lut_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36734\,
            in2 => \N__36728\,
            in3 => \N__48729\,
            lcout => OPEN,
            ltout => \n30_adj_1535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i6_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40198\,
            in1 => \_gnd_net_\,
            in2 => \N__37283\,
            in3 => \N__54077\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57812\,
            ce => \N__42723\,
            sr => \N__42851\
        );

    \ADC_VDC.genclk.i18784_4_lut_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__37276\,
            in1 => \N__37264\,
            in2 => \N__37253\,
            in3 => \N__37231\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n21211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i18825_4_lut_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37085\,
            in1 => \N__37145\,
            in2 => \N__37220\,
            in3 => \N__37019\,
            lcout => \ADC_VDC.genclk.n21205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_adj_25_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37198\,
            in1 => \N__37186\,
            in2 => \N__37175\,
            in3 => \N__37156\,
            lcout => \ADC_VDC.genclk.n26_adj_1408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_adj_24_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37135\,
            in1 => \N__37123\,
            in2 => \N__37112\,
            in3 => \N__37096\,
            lcout => \ADC_VDC.genclk.n28_adj_1407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_adj_26_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__37060\,
            in2 => \N__37049\,
            in3 => \N__37030\,
            lcout => \ADC_VDC.genclk.n27_adj_1409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i0_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37013\,
            in1 => \N__54082\,
            in2 => \_gnd_net_\,
            in3 => \N__50761\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i4_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54080\,
            in1 => \N__40620\,
            in2 => \_gnd_net_\,
            in3 => \N__37001\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i7_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51383\,
            in1 => \N__37403\,
            in2 => \_gnd_net_\,
            in3 => \N__54085\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i6_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54081\,
            in1 => \N__40215\,
            in2 => \_gnd_net_\,
            in3 => \N__37385\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51032\,
            in1 => \N__37370\,
            in2 => \_gnd_net_\,
            in3 => \N__54084\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i3_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54079\,
            in1 => \N__40757\,
            in2 => \_gnd_net_\,
            in3 => \N__37355\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i2_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47221\,
            in1 => \N__37340\,
            in2 => \_gnd_net_\,
            in3 => \N__54083\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \comm_buf_3__i1_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54078\,
            in1 => \N__45362\,
            in2 => \_gnd_net_\,
            in3 => \N__37322\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57820\,
            ce => \N__37304\,
            sr => \N__37292\
        );

    \mux_143_Mux_0_i1_3_lut_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41500\,
            in1 => \N__41157\,
            in2 => \_gnd_net_\,
            in3 => \N__54373\,
            lcout => OPEN,
            ltout => \n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__50680\,
            in1 => \N__37553\,
            in2 => \N__37286\,
            in3 => \N__37526\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57824\,
            ce => \N__46218\,
            sr => \N__46115\
        );

    \i18722_2_lut_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50702\,
            in2 => \_gnd_net_\,
            in3 => \N__54370\,
            lcout => n20970,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_0_i2_3_lut_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54372\,
            in1 => \_gnd_net_\,
            in2 => \N__37571\,
            in3 => \N__37562\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_0_i4_3_lut_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37547\,
            in1 => \N__37457\,
            in2 => \_gnd_net_\,
            in3 => \N__54371\,
            lcout => OPEN,
            ltout => \n4_adj_1507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19366_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__50679\,
            in1 => \N__37535\,
            in2 => \N__37529\,
            in3 => \N__50545\,
            lcout => n21980,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19011_2_lut_3_lut_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__50544\,
            in1 => \N__50678\,
            in2 => \_gnd_net_\,
            in3 => \N__43059\,
            lcout => OPEN,
            ltout => \n21116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010110011"
        )
    port map (
            in0 => \N__54369\,
            in1 => \N__54075\,
            in2 => \N__37520\,
            in3 => \N__37512\,
            lcout => n12_adj_1602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i0_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__54071\,
            in2 => \_gnd_net_\,
            in3 => \N__50777\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i7_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54070\,
            in1 => \_gnd_net_\,
            in2 => \N__51398\,
            in3 => \N__37451\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i6_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40233\,
            in1 => \N__54074\,
            in2 => \_gnd_net_\,
            in3 => \N__37433\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i5_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54069\,
            in1 => \_gnd_net_\,
            in2 => \N__51047\,
            in3 => \N__37421\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i4_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40638\,
            in1 => \N__54073\,
            in2 => \_gnd_net_\,
            in3 => \N__37739\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i3_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54068\,
            in1 => \N__40792\,
            in2 => \_gnd_net_\,
            in3 => \N__37709\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i2_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47234\,
            in1 => \N__54072\,
            in2 => \_gnd_net_\,
            in3 => \N__37688\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \comm_buf_4__i1_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54067\,
            in1 => \N__45363\,
            in2 => \_gnd_net_\,
            in3 => \N__37667\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57833\,
            ce => \N__37646\,
            sr => \N__37634\
        );

    \mux_143_Mux_3_i1_3_lut_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37969\,
            in1 => \N__54331\,
            in2 => \_gnd_net_\,
            in3 => \N__44259\,
            lcout => OPEN,
            ltout => \n1_adj_1589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__37808\,
            in1 => \N__37601\,
            in2 => \N__37622\,
            in3 => \N__50667\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57843\,
            ce => \N__46212\,
            sr => \N__46141\
        );

    \i19059_2_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54329\,
            in2 => \_gnd_net_\,
            in3 => \N__37619\,
            lcout => OPEN,
            ltout => \n21296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__50533\,
            in1 => \N__37577\,
            in2 => \N__37604\,
            in3 => \N__50666\,
            lcout => n22154,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_3_i4_3_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37595\,
            in1 => \N__54328\,
            in2 => \_gnd_net_\,
            in3 => \N__37589\,
            lcout => n4_adj_1591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_3_i2_3_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54330\,
            in1 => \N__37832\,
            in2 => \_gnd_net_\,
            in3 => \N__37823\,
            lcout => n2_adj_1590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18879_3_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54327\,
            in2 => \N__43271\,
            in3 => \N__50532\,
            lcout => OPEN,
            ltout => \n21102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i40_4_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__45193\,
            in1 => \N__54022\,
            in2 => \N__37802\,
            in3 => \N__37799\,
            lcout => n16_adj_1599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_6_i26_3_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56007\,
            in1 => \N__37787\,
            in2 => \_gnd_net_\,
            in3 => \N__46522\,
            lcout => OPEN,
            ltout => \n26_adj_1505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18316_4_lut_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__48153\,
            in1 => \N__37766\,
            in2 => \N__37751\,
            in3 => \N__56008\,
            lcout => OPEN,
            ltout => \n20930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19424_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__37991\,
            in1 => \N__48685\,
            in2 => \N__37748\,
            in3 => \N__48954\,
            lcout => OPEN,
            ltout => \n21962_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21962_bdd_4_lut_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__48686\,
            in1 => \N__38030\,
            in2 => \N__37745\,
            in3 => \N__38324\,
            lcout => OPEN,
            ltout => \n21965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i6_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54086\,
            in1 => \_gnd_net_\,
            in2 => \N__37742\,
            in3 => \N__40244\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57853\,
            ce => \N__47054\,
            sr => \N__46969\
        );

    \mux_135_Mux_6_i19_3_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38108\,
            in1 => \N__38076\,
            in2 => \_gnd_net_\,
            in3 => \N__56006\,
            lcout => OPEN,
            ltout => \n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18340_3_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38051\,
            in2 => \N__38033\,
            in3 => \N__48152\,
            lcout => n20954,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18315_3_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48151\,
            in1 => \_gnd_net_\,
            in2 => \N__38021\,
            in3 => \N__46331\,
            lcout => n20929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40797\,
            in1 => \N__54087\,
            in2 => \_gnd_net_\,
            in3 => \N__37886\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57863\,
            ce => \N__47069\,
            sr => \N__47000\
        );

    \i18270_3_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48312\,
            in1 => \N__47708\,
            in2 => \_gnd_net_\,
            in3 => \N__37931\,
            lcout => OPEN,
            ltout => \n20884_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19557_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__48597\,
            in1 => \N__49075\,
            in2 => \N__37907\,
            in3 => \N__37838\,
            lcout => OPEN,
            ltout => \n22124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22124_bdd_4_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__37904\,
            in1 => \N__38300\,
            in2 => \N__37889\,
            in3 => \N__48598\,
            lcout => n22127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_3_i26_3_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37876\,
            in1 => \N__56269\,
            in2 => \_gnd_net_\,
            in3 => \N__47731\,
            lcout => OPEN,
            ltout => \n26_adj_1514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18271_4_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__56270\,
            in1 => \N__37862\,
            in2 => \N__37841\,
            in3 => \N__48310\,
            lcout => n20885,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18265_3_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38237\,
            in1 => \N__38315\,
            in2 => \_gnd_net_\,
            in3 => \N__48311\,
            lcout => n20879,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_3_i19_3_lut_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__56268\,
            in1 => \N__38286\,
            in2 => \_gnd_net_\,
            in3 => \N__38258\,
            lcout => n19_adj_1513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19533_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__48315\,
            in1 => \N__49050\,
            in2 => \N__52571\,
            in3 => \N__38198\,
            lcout => OPEN,
            ltout => \n22178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22178_bdd_4_lut_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49051\,
            in1 => \N__49283\,
            in2 => \N__38231\,
            in3 => \N__46724\,
            lcout => OPEN,
            ltout => \n22181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1547870_i1_3_lut_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38618\,
            in2 => \N__38228\,
            in3 => \N__48701\,
            lcout => OPEN,
            ltout => \n30_adj_1511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40650\,
            in1 => \_gnd_net_\,
            in2 => \N__38225\,
            in3 => \N__54088\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57873\,
            ce => \N__47071\,
            sr => \N__46995\
        );

    \mux_135_Mux_4_i26_3_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38222\,
            in1 => \N__56184\,
            in2 => \_gnd_net_\,
            in3 => \N__46740\,
            lcout => n26_adj_1510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19400_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000101100"
        )
    port map (
            in0 => \N__38192\,
            in1 => \N__48314\,
            in2 => \N__49127\,
            in3 => \N__38186\,
            lcout => OPEN,
            ltout => \n22010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22010_bdd_4_lut_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49049\,
            in1 => \N__38161\,
            in2 => \N__38126\,
            in3 => \N__38123\,
            lcout => n22013,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_228_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__54764\,
            in1 => \N__49593\,
            in2 => \N__39215\,
            in3 => \N__46585\,
            lcout => n12441,
            ltout => \n12441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__45456\,
            in1 => \N__49630\,
            in2 => \N__38612\,
            in3 => \N__43395\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6464_3_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45454\,
            in1 => \N__38593\,
            in2 => \_gnd_net_\,
            in3 => \N__41746\,
            lcout => n8_adj_1567,
            ltout => \n8_adj_1567_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__54765\,
            in1 => \N__49595\,
            in2 => \N__38609\,
            in3 => \N__42200\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49594\,
            in1 => \N__49344\,
            in2 => \N__46410\,
            in3 => \N__38839\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i1_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__38388\,
            in1 => \N__45457\,
            in2 => \N__38579\,
            in3 => \N__38480\,
            lcout => buf_dds1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15262_2_lut_3_lut_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__54124\,
            in2 => \_gnd_net_\,
            in3 => \N__52434\,
            lcout => n14_adj_1550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i4_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__49592\,
            in1 => \N__44173\,
            in2 => \N__44440\,
            in3 => \N__39016\,
            lcout => \VDC_RNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18339_3_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38359\,
            in1 => \N__38336\,
            in2 => \_gnd_net_\,
            in3 => \N__48313\,
            lcout => n20953,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_239_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110111"
        )
    port map (
            in0 => \N__41748\,
            in1 => \N__54763\,
            in2 => \N__49700\,
            in3 => \N__39157\,
            lcout => n12312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i6_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43154\,
            in1 => \N__44434\,
            in2 => \N__45012\,
            in3 => \N__49590\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_4_i23_3_lut_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39015\,
            in1 => \N__56183\,
            in2 => \_gnd_net_\,
            in3 => \N__38999\,
            lcout => n23_adj_1538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i11_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49591\,
            in1 => \N__40449\,
            in2 => \N__44301\,
            in3 => \N__38968\,
            lcout => buf_dds0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_67_i14_2_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38861\,
            in2 => \_gnd_net_\,
            in3 => \N__38835\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_170_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38813\,
            in1 => \N__49282\,
            in2 => \N__38795\,
            in3 => \N__43396\,
            lcout => n18_adj_1611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i4_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__38741\,
            in1 => \N__54871\,
            in2 => \N__49772\,
            in3 => \N__38725\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_4_i15_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__54870\,
            in1 => \N__38740\,
            in2 => \N__38726\,
            in3 => \N__49682\,
            lcout => \data_index_9_N_216_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_2_i15_4_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54887\,
            in1 => \N__39442\,
            in2 => \N__49771\,
            in3 => \N__39431\,
            lcout => \data_index_9_N_216_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39317\,
            in1 => \N__47413\,
            in2 => \_gnd_net_\,
            in3 => \N__42013\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__49356\,
            in1 => \N__49638\,
            in2 => \N__47795\,
            in3 => \N__46048\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39284\,
            in1 => \N__47414\,
            in2 => \_gnd_net_\,
            in3 => \N__44529\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__39257\,
            in1 => \N__39239\,
            in2 => \N__49181\,
            in3 => \N__46278\,
            lcout => n22_adj_1620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15172_2_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42326\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_193_i9_2_lut_3_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__48359\,
            in1 => \N__56296\,
            in2 => \_gnd_net_\,
            in3 => \N__49099\,
            lcout => n9_adj_1415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41765\,
            in1 => \_gnd_net_\,
            in2 => \N__39200\,
            in3 => \N__47412\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18828_2_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56297\,
            in2 => \_gnd_net_\,
            in3 => \N__41764\,
            lcout => n21048,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44078\,
            in1 => \N__47411\,
            in2 => \_gnd_net_\,
            in3 => \N__42039\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__45566\,
            in1 => \N__44439\,
            in2 => \N__44643\,
            in3 => \N__49776\,
            lcout => \DDS_RNG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_3_lut_3_lut_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__54169\,
            in1 => \N__52407\,
            in2 => \_gnd_net_\,
            in3 => \N__53581\,
            lcout => n10_adj_1613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i0_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42353\,
            in2 => \_gnd_net_\,
            in3 => \N__39473\,
            lcout => dds0_mclkcnt_0,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => n19498,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i1_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42391\,
            in2 => \_gnd_net_\,
            in3 => \N__39470\,
            lcout => dds0_mclkcnt_1,
            ltout => OPEN,
            carryin => n19498,
            carryout => n19499,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i2_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42365\,
            in2 => \_gnd_net_\,
            in3 => \N__39467\,
            lcout => dds0_mclkcnt_2,
            ltout => OPEN,
            carryin => n19499,
            carryout => n19500,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i3_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42416\,
            in2 => \_gnd_net_\,
            in3 => \N__39464\,
            lcout => dds0_mclkcnt_3,
            ltout => OPEN,
            carryin => n19500,
            carryout => n19501,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i4_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42377\,
            in2 => \_gnd_net_\,
            in3 => \N__39461\,
            lcout => dds0_mclkcnt_4,
            ltout => OPEN,
            carryin => n19501,
            carryout => n19502,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i5_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42404\,
            in2 => \_gnd_net_\,
            in3 => \N__39458\,
            lcout => dds0_mclkcnt_5,
            ltout => OPEN,
            carryin => n19502,
            carryout => n19503,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i6_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39455\,
            in2 => \_gnd_net_\,
            in3 => \N__39596\,
            lcout => dds0_mclkcnt_6,
            ltout => OPEN,
            carryin => n19503,
            carryout => n19504,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3783__i7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42338\,
            in2 => \_gnd_net_\,
            in3 => \N__39593\,
            lcout => dds0_mclkcnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclkcnt_i7_3783__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secclk_cnt_3776_3777__i1_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39590\,
            in2 => \_gnd_net_\,
            in3 => \N__39578\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => n19509,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i2_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39574\,
            in2 => \_gnd_net_\,
            in3 => \N__39560\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n19509,
            carryout => n19510,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i3_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39557\,
            in2 => \_gnd_net_\,
            in3 => \N__39545\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n19510,
            carryout => n19511,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i4_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39542\,
            in2 => \_gnd_net_\,
            in3 => \N__39530\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n19511,
            carryout => n19512,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i5_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39527\,
            in2 => \_gnd_net_\,
            in3 => \N__39515\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n19512,
            carryout => n19513,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39512\,
            in2 => \_gnd_net_\,
            in3 => \N__39500\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n19513,
            carryout => n19514,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i7_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39497\,
            in2 => \_gnd_net_\,
            in3 => \N__39485\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n19514,
            carryout => n19515,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i8_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39725\,
            in2 => \_gnd_net_\,
            in3 => \N__39713\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n19515,
            carryout => n19516,
            clk => \N__45084\,
            ce => 'H',
            sr => \N__39763\
        );

    \secclk_cnt_3776_3777__i9_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39710\,
            in2 => \_gnd_net_\,
            in3 => \N__39698\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => n19517,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i10_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39695\,
            in2 => \_gnd_net_\,
            in3 => \N__39683\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n19517,
            carryout => n19518,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i11_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39679\,
            in2 => \_gnd_net_\,
            in3 => \N__39665\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n19518,
            carryout => n19519,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i12_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39662\,
            in2 => \_gnd_net_\,
            in3 => \N__39650\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n19519,
            carryout => n19520,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i13_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39646\,
            in2 => \_gnd_net_\,
            in3 => \N__39632\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n19520,
            carryout => n19521,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i14_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39628\,
            in2 => \_gnd_net_\,
            in3 => \N__39614\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n19521,
            carryout => n19522,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i15_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39611\,
            in2 => \_gnd_net_\,
            in3 => \N__39599\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n19522,
            carryout => n19523,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i16_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39887\,
            in2 => \_gnd_net_\,
            in3 => \N__39875\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n19523,
            carryout => n19524,
            clk => \N__45086\,
            ce => 'H',
            sr => \N__39756\
        );

    \secclk_cnt_3776_3777__i17_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39872\,
            in2 => \_gnd_net_\,
            in3 => \N__39860\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => n19525,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i18_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39857\,
            in2 => \_gnd_net_\,
            in3 => \N__39845\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n19525,
            carryout => n19526,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i19_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39841\,
            in2 => \_gnd_net_\,
            in3 => \N__39827\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n19526,
            carryout => n19527,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i20_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39824\,
            in2 => \_gnd_net_\,
            in3 => \N__39812\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n19527,
            carryout => n19528,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i21_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39809\,
            in2 => \_gnd_net_\,
            in3 => \N__39797\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n19528,
            carryout => n19529,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i22_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39794\,
            in2 => \_gnd_net_\,
            in3 => \N__39782\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n19529,
            carryout => n19530,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \secclk_cnt_3776_3777__i23_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39776\,
            in2 => \_gnd_net_\,
            in3 => \N__39779\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45090\,
            ce => 'H',
            sr => \N__39764\
        );

    \comm_spi.data_rx_i3_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42605\,
            in1 => \N__47181\,
            in2 => \_gnd_net_\,
            in3 => \N__40523\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i4_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__40520\,
            in1 => \N__40736\,
            in2 => \_gnd_net_\,
            in3 => \N__42606\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i5_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42607\,
            in1 => \N__40599\,
            in2 => \_gnd_net_\,
            in3 => \N__40524\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i6_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__40521\,
            in1 => \N__50994\,
            in2 => \_gnd_net_\,
            in3 => \N__42608\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i7_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42609\,
            in1 => \N__40197\,
            in2 => \_gnd_net_\,
            in3 => \N__40525\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i2_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__40519\,
            in1 => \N__45321\,
            in2 => \_gnd_net_\,
            in3 => \N__42604\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \comm_spi.data_rx_i1_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__42603\,
            in1 => \N__40522\,
            in2 => \_gnd_net_\,
            in3 => \N__50775\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57050\,
            ce => 'H',
            sr => \N__56858\
        );

    \ADC_VDC.genclk.t_clk_24_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40175\,
            lcout => \VDC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t_clk_24C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__42535\,
            in1 => \N__42557\,
            in2 => \_gnd_net_\,
            in3 => \N__42573\,
            lcout => \comm_spi.n16869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12402_3_lut_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__40570\,
            in1 => \N__46219\,
            in2 => \_gnd_net_\,
            in3 => \N__54528\,
            lcout => n14815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18892_3_lut_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__54055\,
            in1 => \N__41102\,
            in2 => \_gnd_net_\,
            in3 => \N__40571\,
            lcout => OPEN,
            ltout => \n21506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18269_4_lut_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__43217\,
            in1 => \N__45644\,
            in2 => \N__40424\,
            in3 => \N__52326\,
            lcout => n20883,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12353_2_lut_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__54529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42689\,
            lcout => n14766,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22028_bdd_4_lut_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__40421\,
            in1 => \N__40388\,
            in2 => \N__40406\,
            in3 => \N__49077\,
            lcout => n22031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19429_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__48316\,
            in1 => \N__45233\,
            in2 => \N__40925\,
            in3 => \N__49076\,
            lcout => n22028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19459_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56368\,
            in1 => \N__41323\,
            in2 => \N__40381\,
            in3 => \N__48317\,
            lcout => OPEN,
            ltout => \n22088_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22088_bdd_4_lut_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48318\,
            in1 => \N__40340\,
            in2 => \N__40307\,
            in3 => \N__40304\,
            lcout => OPEN,
            ltout => \n22091_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18230_3_lut_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49078\,
            in1 => \_gnd_net_\,
            in2 => \N__40274\,
            in3 => \N__40271\,
            lcout => OPEN,
            ltout => \n20844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1543649_i1_3_lut_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40256\,
            in2 => \N__40250\,
            in3 => \N__48742\,
            lcout => OPEN,
            ltout => \n30_adj_1539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i4_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40619\,
            in1 => \_gnd_net_\,
            in2 => \N__40574\,
            in3 => \N__54036\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57825\,
            ce => \N__42717\,
            sr => \N__42831\
        );

    \i1_2_lut_3_lut_4_lut_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__51828\,
            in1 => \N__50669\,
            in2 => \N__51669\,
            in3 => \N__40562\,
            lcout => n20596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_68_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40563\,
            in1 => \N__53549\,
            in2 => \N__51843\,
            in3 => \N__51642\,
            lcout => n20621,
            ltout => \n20621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_248_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40535\,
            in3 => \N__50538\,
            lcout => OPEN,
            ltout => \n25_adj_1619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_231_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__50670\,
            in1 => \N__54352\,
            in2 => \N__40532\,
            in3 => \N__54030\,
            lcout => n4_adj_1616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__40529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42617\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__56854\
        );

    \i22_4_lut_4_lut_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000100010"
        )
    port map (
            in0 => \N__53519\,
            in1 => \N__54031\,
            in2 => \N__51844\,
            in3 => \N__51646\,
            lcout => n7_adj_1609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110011"
        )
    port map (
            in0 => \N__53520\,
            in1 => \N__54032\,
            in2 => \N__51845\,
            in3 => \N__51647\,
            lcout => n20717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22082_bdd_4_lut_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48293\,
            in1 => \N__40484\,
            in2 => \N__40456\,
            in3 => \N__40871\,
            lcout => n22085,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19449_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56185\,
            in1 => \N__41077\,
            in2 => \N__40909\,
            in3 => \N__48292\,
            lcout => n22082,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_3_i26_3_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40865\,
            in1 => \N__56186\,
            in2 => \_gnd_net_\,
            in3 => \N__41786\,
            lcout => OPEN,
            ltout => \n26_adj_1541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18223_4_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__56187\,
            in1 => \N__40844\,
            in2 => \N__40829\,
            in3 => \N__48294\,
            lcout => OPEN,
            ltout => \n20837_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19464_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__44501\,
            in1 => \N__48736\,
            in2 => \N__40826\,
            in3 => \N__49053\,
            lcout => OPEN,
            ltout => \n22094_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22094_bdd_4_lut_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__48737\,
            in1 => \N__40823\,
            in2 => \N__40817\,
            in3 => \N__40814\,
            lcout => OPEN,
            ltout => \n22097_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i3_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40758\,
            in2 => \N__40700\,
            in3 => \N__53994\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57844\,
            ce => \N__42724\,
            sr => \N__42852\
        );

    \i6988_2_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__52390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54006\,
            lcout => n9321,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_217_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__54637\,
            in1 => \N__51542\,
            in2 => \N__51605\,
            in3 => \N__52393\,
            lcout => n11406,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \flagcntwd_313_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54008\,
            in2 => \_gnd_net_\,
            in3 => \N__53504\,
            lcout => flagcntwd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57854\,
            ce => \N__40667\,
            sr => \N__51212\
        );

    \i1_2_lut_3_lut_adj_301_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__52391\,
            in1 => \N__54007\,
            in2 => \_gnd_net_\,
            in3 => \N__54635\,
            lcout => n12242,
            ltout => \n12242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_86_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__54636\,
            in1 => \_gnd_net_\,
            in2 => \N__41108\,
            in3 => \N__52392\,
            lcout => n20599,
            ltout => \n20599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_236_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__50925\,
            in1 => \N__53503\,
            in2 => \N__41105\,
            in3 => \N__43238\,
            lcout => n12047,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_254_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__47911\,
            in1 => \N__50552\,
            in2 => \_gnd_net_\,
            in3 => \N__47866\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49449\,
            in1 => \N__41390\,
            in2 => \N__44302\,
            in3 => \N__41073\,
            lcout => \IAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12241_2_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__41053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41885\,
            lcout => n14663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12360_2_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54654\,
            in2 => \_gnd_net_\,
            in3 => \N__47029\,
            lcout => n14773,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18728_2_lut_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40958\,
            in2 => \_gnd_net_\,
            in3 => \N__56324\,
            lcout => n20973,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18739_2_lut_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40946\,
            lcout => n20983,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41389\,
            in1 => \N__44127\,
            in2 => \N__49833\,
            in3 => \N__41322\,
            lcout => \VAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18816_2_lut_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__56322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47510\,
            lcout => n21046,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21998_bdd_4_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__41204\,
            in1 => \N__41291\,
            in2 => \N__46469\,
            in3 => \N__49106\,
            lcout => n22001,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19385_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__49105\,
            in1 => \N__41270\,
            in2 => \N__41258\,
            in3 => \N__48337\,
            lcout => n22004,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_0_i26_3_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41233\,
            in1 => \N__56271\,
            in2 => \_gnd_net_\,
            in3 => \N__46492\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19380_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__49104\,
            in1 => \N__41216\,
            in2 => \N__41207\,
            in3 => \N__48336\,
            lcout => n21998,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22004_bdd_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__41198\,
            in1 => \N__41186\,
            in2 => \N__52157\,
            in3 => \N__49107\,
            lcout => OPEN,
            ltout => \n22007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1548473_i1_3_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48607\,
            in2 => \N__41180\,
            in3 => \N__41177\,
            lcout => OPEN,
            ltout => \n30_adj_1486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i0_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54051\,
            in2 => \N__41171\,
            in3 => \N__50771\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57874\,
            ce => \N__47053\,
            sr => \N__46970\
        );

    \n21992_bdd_4_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__41591\,
            in1 => \N__41657\,
            in2 => \N__48423\,
            in3 => \N__49979\,
            lcout => n21995,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19390_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__56319\,
            in1 => \N__41630\,
            in2 => \N__48365\,
            in3 => \N__43901\,
            lcout => n21992,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18303_3_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41585\,
            in1 => \N__56320\,
            in2 => \_gnd_net_\,
            in3 => \N__43460\,
            lcout => OPEN,
            ltout => \n20917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18305_4_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__56321\,
            in1 => \N__41564\,
            in2 => \N__41555\,
            in3 => \N__48408\,
            lcout => OPEN,
            ltout => \n20919_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19567_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__49013\,
            in1 => \N__41552\,
            in2 => \N__41546\,
            in3 => \N__48700\,
            lcout => OPEN,
            ltout => \n22220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22220_bdd_4_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__41543\,
            in1 => \N__41531\,
            in2 => \N__41516\,
            in3 => \N__48688\,
            lcout => OPEN,
            ltout => \n22223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54052\,
            in2 => \N__41513\,
            in3 => \N__50782\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57887\,
            ce => \N__42722\,
            sr => \N__42857\
        );

    \i19053_4_lut_4_lut_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101101011"
        )
    port map (
            in0 => \N__56318\,
            in1 => \N__48687\,
            in2 => \N__48364\,
            in3 => \N__49012\,
            lcout => n21094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46491\,
            in2 => \N__41441\,
            in3 => \_gnd_net_\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => n19354,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46767\,
            in2 => \_gnd_net_\,
            in3 => \N__41684\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n19354,
            carryout => n19355,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46845\,
            in2 => \_gnd_net_\,
            in3 => \N__41681\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n19355,
            carryout => n19356,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47730\,
            in2 => \_gnd_net_\,
            in3 => \N__41678\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n19356,
            carryout => n19357,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46744\,
            in2 => \_gnd_net_\,
            in3 => \N__41675\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n19357,
            carryout => n19358,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i5_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47753\,
            in2 => \_gnd_net_\,
            in3 => \N__41672\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n19358,
            carryout => n19359,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i6_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46521\,
            in2 => \_gnd_net_\,
            in3 => \N__41669\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n19359,
            carryout => n19360,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i7_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49225\,
            in2 => \_gnd_net_\,
            in3 => \N__41666\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n19360,
            carryout => n19361,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__41887\,
            sr => \N__41832\
        );

    \data_cntvec_i0_i8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43459\,
            in2 => \_gnd_net_\,
            in3 => \N__41663\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => n19362,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i9_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47530\,
            in2 => \_gnd_net_\,
            in3 => \N__41660\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n19362,
            carryout => n19363,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i10_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42061\,
            in2 => \_gnd_net_\,
            in3 => \N__41906\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n19363,
            carryout => n19364,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i11_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41785\,
            in2 => \_gnd_net_\,
            in3 => \N__41903\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n19364,
            carryout => n19365,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i12_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42080\,
            in2 => \_gnd_net_\,
            in3 => \N__41900\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n19365,
            carryout => n19366,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i13_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43438\,
            in2 => \_gnd_net_\,
            in3 => \N__41897\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n19366,
            carryout => n19367,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i14_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41798\,
            in2 => \_gnd_net_\,
            in3 => \N__41894\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n19367,
            carryout => n19368,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \data_cntvec_i0_i15_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47485\,
            in2 => \_gnd_net_\,
            in3 => \N__41891\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__41888\,
            sr => \N__41828\
        );

    \i7_4_lut_adj_182_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__41784\,
            in2 => \N__44536\,
            in3 => \N__41763\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6414_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52489\,
            in1 => \N__41949\,
            in2 => \_gnd_net_\,
            in3 => \N__41750\,
            lcout => n8_adj_1559,
            ltout => \n8_adj_1559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_6_i15_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__41983\,
            in1 => \N__54868\,
            in2 => \N__42305\,
            in3 => \N__49521\,
            lcout => \data_index_9_N_216_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_365_Mux_1_i15_4_lut_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54867\,
            in1 => \N__42212\,
            in2 => \N__49629\,
            in3 => \N__42199\,
            lcout => \data_index_9_N_216_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__47135\,
            in1 => \N__49366\,
            in2 => \N__46288\,
            in3 => \N__49522\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_184_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__42079\,
            in1 => \N__42060\,
            in2 => \N__42040\,
            in3 => \N__42009\,
            lcout => n21_adj_1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__41993\,
            in1 => \N__54869\,
            in2 => \N__41987\,
            in3 => \N__49523\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__56852\,
            in1 => \N__55311\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_771\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_cnt_3772_3773__i1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42512\,
            in2 => \_gnd_net_\,
            in3 => \N__41915\,
            lcout => clk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => n19505,
            clk => \N__45083\,
            ce => 'H',
            sr => \N__43838\
        );

    \clk_cnt_3772_3773__i2_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42487\,
            in2 => \_gnd_net_\,
            in3 => \N__41912\,
            lcout => clk_cnt_1,
            ltout => OPEN,
            carryin => n19505,
            carryout => n19506,
            clk => \N__45083\,
            ce => 'H',
            sr => \N__43838\
        );

    \clk_cnt_3772_3773__i3_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42457\,
            in2 => \_gnd_net_\,
            in3 => \N__41909\,
            lcout => clk_cnt_2,
            ltout => OPEN,
            carryin => n19506,
            carryout => n19507,
            clk => \N__45083\,
            ce => 'H',
            sr => \N__43838\
        );

    \clk_cnt_3772_3773__i4_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42473\,
            in2 => \_gnd_net_\,
            in3 => \N__42518\,
            lcout => clk_cnt_3,
            ltout => OPEN,
            carryin => n19507,
            carryout => n19508,
            clk => \N__45083\,
            ce => 'H',
            sr => \N__43838\
        );

    \clk_cnt_3772_3773__i5_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42500\,
            in2 => \_gnd_net_\,
            in3 => \N__42515\,
            lcout => clk_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45083\,
            ce => 'H',
            sr => \N__43838\
        );

    \i1_2_lut_adj_232_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42499\,
            lcout => OPEN,
            ltout => \n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_234_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42488\,
            in1 => \N__42472\,
            in2 => \N__42461\,
            in3 => \N__42458\,
            lcout => n14730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_3_i23_3_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44197\,
            in1 => \N__56334\,
            in2 => \_gnd_net_\,
            in3 => \N__42443\,
            lcout => n23_adj_1540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42415\,
            in1 => \N__42403\,
            in2 => \N__42392\,
            in3 => \N__42376\,
            lcout => OPEN,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_165_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42364\,
            in1 => \N__42352\,
            in2 => \N__42341\,
            in3 => \N__42337\,
            lcout => n20543,
            ltout => \n20543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclk_304_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45028\,
            in2 => \N__42320\,
            in3 => \N__42317\,
            lcout => dds0_mclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclk_304C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__44753\,
            in1 => \N__44845\,
            in2 => \N__44870\,
            in3 => \N__44828\,
            lcout => \SIG_DDS.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57960\,
            ce => \N__50176\,
            sr => \N__44765\
        );

    \SIG_DDS.bit_cnt_i1_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44862\,
            in2 => \_gnd_net_\,
            in3 => \N__44751\,
            lcout => \SIG_DDS.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57960\,
            ce => \N__50176\,
            sr => \N__44765\
        );

    \SIG_DDS.bit_cnt_i2_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44752\,
            in1 => \_gnd_net_\,
            in2 => \N__44869\,
            in3 => \N__44844\,
            lcout => \SIG_DDS.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57960\,
            ce => \N__50176\,
            sr => \N__44765\
        );

    \SIG_DDS.dds_state_i2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50233\,
            in2 => \_gnd_net_\,
            in3 => \N__50156\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18840_2_lut_LC_16_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42638\,
            in2 => \_gnd_net_\,
            in3 => \N__56370\,
            lcout => n21038,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_3778__i3_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__42575\,
            in1 => \N__42610\,
            in2 => \N__42542\,
            in3 => \N__42560\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3778__i3C_net\,
            ce => 'H',
            sr => \N__56823\
        );

    \comm_spi.bit_cnt_3778__i2_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__42559\,
            in1 => \N__42538\,
            in2 => \_gnd_net_\,
            in3 => \N__42574\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3778__i3C_net\,
            ce => 'H',
            sr => \N__56823\
        );

    \comm_spi.bit_cnt_3778__i1_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42558\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3778__i3C_net\,
            ce => 'H',
            sr => \N__56823\
        );

    \comm_spi.bit_cnt_3778__i0_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42536\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3778__i3C_net\,
            ce => 'H',
            sr => \N__56823\
        );

    \comm_buf_0__i7_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51342\,
            in1 => \N__54035\,
            in2 => \_gnd_net_\,
            in3 => \N__42893\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57826\,
            ce => \N__42721\,
            sr => \N__42847\
        );

    \comm_buf_0__i5_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54033\,
            in1 => \N__50995\,
            in2 => \_gnd_net_\,
            in3 => \N__42878\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57826\,
            ce => \N__42721\,
            sr => \N__42847\
        );

    \comm_buf_0__i1_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45322\,
            in1 => \N__54034\,
            in2 => \_gnd_net_\,
            in3 => \N__44003\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57826\,
            ce => \N__42721\,
            sr => \N__42847\
        );

    \i18822_2_lut_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45742\,
            in2 => \_gnd_net_\,
            in3 => \N__53518\,
            lcout => OPEN,
            ltout => \n21199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001010101"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__49626\,
            in2 => \N__42791\,
            in3 => \N__54559\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57835\,
            ce => \N__45749\,
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__54029\,
            in1 => \N__50885\,
            in2 => \N__45205\,
            in3 => \N__53516\,
            lcout => n11869,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_105_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52259\,
            in2 => \_gnd_net_\,
            in3 => \N__54558\,
            lcout => n20681,
            ltout => \n20681_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_129_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__45201\,
            in1 => \N__53862\,
            in2 => \N__42788\,
            in3 => \N__53517\,
            lcout => OPEN,
            ltout => \n12108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_233_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__50886\,
            in1 => \N__42778\,
            in2 => \N__42734\,
            in3 => \N__42731\,
            lcout => n11977,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_6_i2_3_lut_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54344\,
            in1 => \N__42659\,
            in2 => \_gnd_net_\,
            in3 => \N__42647\,
            lcout => n2_adj_1584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19041_2_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43205\,
            in2 => \_gnd_net_\,
            in3 => \N__54345\,
            lcout => OPEN,
            ltout => \n21329_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19489_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__50547\,
            in1 => \N__54191\,
            in2 => \N__43187\,
            in3 => \N__50682\,
            lcout => OPEN,
            ltout => \n21986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50683\,
            in1 => \N__43079\,
            in2 => \N__43184\,
            in3 => \N__43181\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57845\,
            ce => \N__46213\,
            sr => \N__46116\
        );

    \mux_143_Mux_6_i1_3_lut_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43136\,
            in1 => \N__52505\,
            in2 => \_gnd_net_\,
            in3 => \N__54343\,
            lcout => n1_adj_1583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_295_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__50546\,
            in1 => \N__43063\,
            in2 => \_gnd_net_\,
            in3 => \N__50681\,
            lcout => OPEN,
            ltout => \n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_156_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__45764\,
            in1 => \N__51568\,
            in2 => \N__43043\,
            in3 => \N__54530\,
            lcout => n12244,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19419_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__54270\,
            in1 => \N__43040\,
            in2 => \N__43025\,
            in3 => \N__50482\,
            lcout => OPEN,
            ltout => \n22046_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22046_bdd_4_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50483\,
            in1 => \N__42972\,
            in2 => \N__42896\,
            in3 => \N__47134\,
            lcout => n22049,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_2_i4_3_lut_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54271\,
            in1 => \N__43328\,
            in2 => \_gnd_net_\,
            in3 => \N__43316\,
            lcout => OPEN,
            ltout => \n4_adj_1593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18187_4_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__50484\,
            in1 => \N__43307\,
            in2 => \N__43283\,
            in3 => \N__54272\,
            lcout => OPEN,
            ltout => \n20801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43280\,
            in2 => \N__43274\,
            in3 => \N__50636\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57855\,
            ce => \N__46205\,
            sr => \N__46133\
        );

    \i18878_3_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__50481\,
            in1 => \N__54269\,
            in2 => \_gnd_net_\,
            in3 => \N__43264\,
            lcout => OPEN,
            ltout => \n21092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i45_4_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__43253\,
            in1 => \N__45194\,
            in2 => \N__43241\,
            in3 => \N__53917\,
            lcout => n20_adj_1610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__49448\,
            in1 => \N__43232\,
            in2 => \_gnd_net_\,
            in3 => \N__54705\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57865\,
            ce => \N__45671\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_308_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53770\,
            in2 => \_gnd_net_\,
            in3 => \N__53495\,
            lcout => OPEN,
            ltout => \n20695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_292_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50906\,
            in1 => \N__51827\,
            in2 => \N__43220\,
            in3 => \N__51670\,
            lcout => n20697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18267_3_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__51825\,
            in1 => \N__53771\,
            in2 => \_gnd_net_\,
            in3 => \N__53496\,
            lcout => n20881,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__53497\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51826\,
            lcout => n14545,
            ltout => \n14545_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_306_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__51671\,
            in1 => \N__53772\,
            in2 => \N__43424\,
            in3 => \N__50907\,
            lcout => n11420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__51394\,
            in1 => \N__54026\,
            in2 => \_gnd_net_\,
            in3 => \N__43850\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57875\,
            ce => \N__47061\,
            sr => \N__46989\
        );

    \mux_135_Mux_1_i26_3_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43420\,
            in1 => \N__56329\,
            in2 => \_gnd_net_\,
            in3 => \N__46768\,
            lcout => OPEN,
            ltout => \n26_adj_1522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19547_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__45839\,
            in1 => \N__48339\,
            in2 => \N__43403\,
            in3 => \N__49114\,
            lcout => OPEN,
            ltout => \n22190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22190_bdd_4_lut_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__43400\,
            in1 => \N__49115\,
            in2 => \N__43376\,
            in3 => \N__46694\,
            lcout => OPEN,
            ltout => \n22193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1546061_i1_3_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43607\,
            in2 => \N__43373\,
            in3 => \N__48727\,
            lcout => OPEN,
            ltout => \n30_adj_1523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i1_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45372\,
            in2 => \N__43370\,
            in3 => \N__54053\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57888\,
            ce => \N__47070\,
            sr => \N__46993\
        );

    \comm_cmd_1__bdd_4_lut_19434_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__43367\,
            in1 => \N__48338\,
            in2 => \N__43352\,
            in3 => \N__49112\,
            lcout => OPEN,
            ltout => \n22064_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22064_bdd_4_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49113\,
            in1 => \N__52609\,
            in2 => \N__43625\,
            in3 => \N__43622\,
            lcout => n22067,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19499_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010110000"
        )
    port map (
            in0 => \N__43601\,
            in1 => \N__49109\,
            in2 => \N__48425\,
            in3 => \N__46619\,
            lcout => OPEN,
            ltout => \n22142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22142_bdd_4_lut_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49110\,
            in1 => \N__43583\,
            in2 => \N__43547\,
            in3 => \N__43544\,
            lcout => n22145,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22130_bdd_4_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__43466\,
            in1 => \N__49111\,
            in2 => \N__47291\,
            in3 => \N__43529\,
            lcout => OPEN,
            ltout => \n22133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1549076_i1_3_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43502\,
            in2 => \N__43496\,
            in3 => \N__48702\,
            lcout => OPEN,
            ltout => \n30_adj_1499_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51054\,
            in2 => \N__43493\,
            in3 => \N__54054\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57900\,
            ce => \N__47068\,
            sr => \N__46994\
        );

    \mux_135_Mux_5_i26_3_lut_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43490\,
            in1 => \N__56325\,
            in2 => \_gnd_net_\,
            in3 => \N__47745\,
            lcout => OPEN,
            ltout => \n26_adj_1498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19494_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__52541\,
            in1 => \N__48295\,
            in2 => \N__43469\,
            in3 => \N__49108\,
            lcout => n22130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_189_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__43458\,
            in1 => \N__47547\,
            in2 => \N__43439\,
            in3 => \N__43899\,
            lcout => OPEN,
            ltout => \n19_adj_1597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_adj_194_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46445\,
            in1 => \N__47687\,
            in2 => \N__43931\,
            in3 => \N__46676\,
            lcout => OPEN,
            ltout => \n29_adj_1635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_196_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44897\,
            in2 => \N__43928\,
            in3 => \N__44354\,
            lcout => n16_adj_1623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__43900\,
            in1 => \_gnd_net_\,
            in2 => \N__44489\,
            in3 => \N__47397\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_339_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44898\,
            in1 => \N__45536\,
            in2 => \_gnd_net_\,
            in3 => \N__43886\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47396\,
            in1 => \N__51118\,
            in2 => \_gnd_net_\,
            in3 => \N__46716\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44050\,
            in1 => \N__47395\,
            in2 => \_gnd_net_\,
            in3 => \N__46310\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57917\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22058_bdd_4_lut_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__43862\,
            in1 => \N__48735\,
            in2 => \N__44921\,
            in3 => \N__49187\,
            lcout => n22061,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_RTD_297_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__43656\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43837\,
            lcout => \clk_RTD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__45080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_181_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__46849\,
            in1 => \N__49224\,
            in2 => \N__49157\,
            in3 => \N__46308\,
            lcout => OPEN,
            ltout => \n22_adj_1568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_192_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44369\,
            in1 => \N__44363\,
            in2 => \N__44357\,
            in3 => \N__47468\,
            lcout => n30_adj_1641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18198_3_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56335\,
            in1 => \N__44348\,
            in2 => \_gnd_net_\,
            in3 => \N__47526\,
            lcout => OPEN,
            ltout => \n20812_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18200_4_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__44327\,
            in1 => \N__48285\,
            in2 => \N__44312\,
            in3 => \N__56336\,
            lcout => n20814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i3_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49739\,
            in1 => \N__44441\,
            in2 => \N__44303\,
            in3 => \N__44193\,
            lcout => \SELIRNG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15254_2_lut_3_lut_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54129\,
            in1 => \N__44139\,
            in2 => \_gnd_net_\,
            in3 => \N__52409\,
            lcout => n14_adj_1571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15261_2_lut_3_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52408\,
            in1 => \N__47133\,
            in2 => \_gnd_net_\,
            in3 => \N__54128\,
            lcout => n14_adj_1549,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__49124\,
            in1 => \N__44594\,
            in2 => \N__48743\,
            in3 => \N__44024\,
            lcout => OPEN,
            ltout => \n22232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22232_bdd_4_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__44018\,
            in1 => \N__44666\,
            in2 => \N__44006\,
            in3 => \N__48734\,
            lcout => n22235,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22226_bdd_4_lut_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__48384\,
            in1 => \N__43991\,
            in2 => \N__43960\,
            in3 => \N__44681\,
            lcout => n22229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22034_bdd_4_lut_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010011000"
        )
    port map (
            in0 => \N__44879\,
            in1 => \N__48370\,
            in2 => \N__44653\,
            in3 => \N__44615\,
            lcout => n22037,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_7_i16_3_lut_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44587\,
            in1 => \N__44563\,
            in2 => \_gnd_net_\,
            in3 => \N__56331\,
            lcout => n16_adj_1503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18222_4_lut_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56332\,
            in1 => \N__48371\,
            in2 => \N__44540\,
            in3 => \N__44507\,
            lcout => n20836,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i0_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44488\,
            in1 => \N__44438\,
            in2 => \_gnd_net_\,
            in3 => \N__49971\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18970_2_lut_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48372\,
            lcout => OPEN,
            ltout => \n21073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18852_4_lut_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__49125\,
            in1 => \N__54736\,
            in2 => \N__44375\,
            in3 => \N__48740\,
            lcout => OPEN,
            ltout => \n21072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__56333\,
            in1 => \N__51442\,
            in2 => \N__44372\,
            in3 => \N__47888\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19135_4_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__50083\,
            in1 => \N__44816\,
            in2 => \N__50362\,
            in3 => \N__50261\,
            lcout => \SIG_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i12483_3_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__50260\,
            in1 => \N__50349\,
            in2 => \_gnd_net_\,
            in3 => \N__50082\,
            lcout => n14900,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_16MHz_I_0_3_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45098\,
            in1 => \N__45032\,
            in2 => \_gnd_net_\,
            in3 => \N__45016\,
            lcout => \DDS_MCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18183_3_lut_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44963\,
            in1 => \N__44927\,
            in2 => \_gnd_net_\,
            in3 => \N__48369\,
            lcout => n20797,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19410_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__56330\,
            in1 => \N__44906\,
            in2 => \N__48409\,
            in3 => \N__47432\,
            lcout => n22034,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i4_4_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44861\,
            in1 => \N__44749\,
            in2 => \N__44846\,
            in3 => \N__50353\,
            lcout => \SIG_DDS.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i18809_2_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44827\,
            in2 => \_gnd_net_\,
            in3 => \N__50223\,
            lcout => \SIG_DDS.n21331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i23_4_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011011"
        )
    port map (
            in0 => \N__50354\,
            in1 => \N__50224\,
            in2 => \N__44815\,
            in3 => \N__50084\,
            lcout => \SIG_DDS.n9_adj_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i0_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__50086\,
            in1 => \N__44750\,
            in2 => \_gnd_net_\,
            in3 => \N__44764\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.MOSI_31_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50085\,
            in1 => \N__44732\,
            in2 => \_gnd_net_\,
            in3 => \N__44692\,
            lcout => \DDS_MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.CS_28_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__50254\,
            in1 => \N__50360\,
            in2 => \_gnd_net_\,
            in3 => \N__50130\,
            lcout => \DDS_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57973\,
            ce => \N__45260\,
            sr => \_gnd_net_\
        );

    \i18846_2_lut_LC_17_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45245\,
            in2 => \_gnd_net_\,
            in3 => \N__56369\,
            lcout => n20984,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_353_Mux_3_i7_4_lut_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__45643\,
            in1 => \N__45799\,
            in2 => \N__45215\,
            in3 => \N__52305\,
            lcout => n17738,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11728_2_lut_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__53957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53563\,
            lcout => n14146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i32_4_lut_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__50855\,
            in1 => \N__53959\,
            in2 => \N__45206\,
            in3 => \N__52306\,
            lcout => OPEN,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__49934\,
            in1 => \N__45134\,
            in2 => \N__45137\,
            in3 => \N__53565\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57836\,
            ce => \N__50813\,
            sr => \N__54836\
        );

    \i33_3_lut_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53564\,
            in1 => \N__45800\,
            in2 => \_gnd_net_\,
            in3 => \N__53958\,
            lcout => n12_adj_1649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_1_i4_3_lut_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45128\,
            in1 => \N__45116\,
            in2 => \_gnd_net_\,
            in3 => \N__54346\,
            lcout => OPEN,
            ltout => \n4_adj_1595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18193_4_lut_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__54347\,
            in1 => \N__45289\,
            in2 => \N__45101\,
            in3 => \N__50534\,
            lcout => n20807,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__45605\,
            in1 => \N__50535\,
            in2 => \N__54374\,
            in3 => \N__45593\,
            lcout => OPEN,
            ltout => \n22052_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22052_bdd_4_lut_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50536\,
            in1 => \N__45537\,
            in2 => \N__45470\,
            in3 => \N__45453\,
            lcout => OPEN,
            ltout => \n22055_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45413\,
            in2 => \N__45407\,
            in3 => \N__50665\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57846\,
            ce => \N__46214\,
            sr => \N__46132\
        );

    \i15005_3_lut_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50663\,
            in1 => \N__45404\,
            in2 => \_gnd_net_\,
            in3 => \N__45912\,
            lcout => OPEN,
            ltout => \n17404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18337_4_lut_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__45392\,
            in1 => \N__50537\,
            in2 => \N__45383\,
            in3 => \N__50664\,
            lcout => OPEN,
            ltout => \n20951_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54351\,
            in2 => \N__45380\,
            in3 => \N__45704\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57846\,
            ce => \N__46214\,
            sr => \N__46132\
        );

    \comm_buf_6__i1_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__51284\,
            in1 => \N__45290\,
            in2 => \N__45376\,
            in3 => \N__54537\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_307_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110101"
        )
    port map (
            in0 => \N__53812\,
            in1 => \N__53537\,
            in2 => \N__51782\,
            in3 => \N__51673\,
            lcout => OPEN,
            ltout => \n4_adj_1598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_84_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__51482\,
            in1 => \N__50834\,
            in2 => \N__45752\,
            in3 => \N__45698\,
            lcout => n20573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i235_2_lut_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__51766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51672\,
            lcout => n1272,
            ltout => \n1272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_353_Mux_1_i8_3_lut_4_lut_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__53538\,
            in1 => \N__45743\,
            in2 => \N__45719\,
            in3 => \N__53813\,
            lcout => n8_adj_1576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22172_bdd_4_lut_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__50414\,
            in1 => \N__45716\,
            in2 => \N__50555\,
            in3 => \N__46355\,
            lcout => n22175,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_299_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__50942\,
            in1 => \N__51476\,
            in2 => \N__51838\,
            in3 => \N__45806\,
            lcout => n20551,
            ltout => \n20551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__51477\,
            in1 => \N__45692\,
            in2 => \N__45683\,
            in3 => \N__45680\,
            lcout => n20575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_1__bdd_4_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__45659\,
            in1 => \N__53921\,
            in2 => \N__45636\,
            in3 => \N__52376\,
            lcout => n22238,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_353_Mux_1_i2_3_lut_4_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__53466\,
            in1 => \N__51839\,
            in2 => \N__54056\,
            in3 => \N__45821\,
            lcout => OPEN,
            ltout => \n2_adj_1575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22238_bdd_4_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__45614\,
            in1 => \N__52377\,
            in2 => \N__45608\,
            in3 => \N__53467\,
            lcout => OPEN,
            ltout => \n22241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i1_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49627\,
            in1 => \N__54722\,
            in2 => \N__45830\,
            in3 => \N__45827\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57866\,
            ce => \N__50951\,
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_296_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__53465\,
            in1 => \N__45820\,
            in2 => \N__51573\,
            in3 => \N__45812\,
            lcout => n4_adj_1614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_309_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111111"
        )
    port map (
            in0 => \N__50493\,
            in1 => \N__47867\,
            in2 => \N__47915\,
            in3 => \N__53774\,
            lcout => n20668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__51692\,
            in1 => \N__51842\,
            in2 => \N__54367\,
            in3 => \N__50495\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57876\,
            ce => \N__45788\,
            sr => \N__45770\
        );

    \comm_index_i0_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__51841\,
            in1 => \N__54320\,
            in2 => \_gnd_net_\,
            in3 => \N__51691\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57876\,
            ce => \N__45788\,
            sr => \N__45770\
        );

    \i1_4_lut_adj_226_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__54707\,
            in1 => \N__53350\,
            in2 => \N__52406\,
            in3 => \N__51550\,
            lcout => n14753,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i2_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__54319\,
            in1 => \N__50494\,
            in2 => \N__50668\,
            in3 => \N__50854\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57876\,
            ce => \N__45788\,
            sr => \N__45770\
        );

    \i3_3_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__52349\,
            in1 => \N__54318\,
            in2 => \_gnd_net_\,
            in3 => \N__53773\,
            lcout => n8_adj_1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_252_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__51549\,
            in1 => \N__52348\,
            in2 => \N__53351\,
            in3 => \N__54706\,
            lcout => n11503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_7_i2_3_lut_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46253\,
            in1 => \N__46241\,
            in2 => \_gnd_net_\,
            in3 => \N__54290\,
            lcout => OPEN,
            ltout => \n2_adj_1581_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__45923\,
            in1 => \N__45965\,
            in2 => \N__46226\,
            in3 => \N__50632\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57889\,
            ce => \N__46198\,
            sr => \N__46142\
        );

    \i18720_2_lut_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51265\,
            in2 => \_gnd_net_\,
            in3 => \N__54287\,
            lcout => n20966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_7_i1_3_lut_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54289\,
            in1 => \N__47630\,
            in2 => \_gnd_net_\,
            in3 => \N__46041\,
            lcout => n1_adj_1580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_143_Mux_7_i4_3_lut_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45959\,
            in1 => \N__45944\,
            in2 => \_gnd_net_\,
            in3 => \N__54288\,
            lcout => OPEN,
            ltout => \n4_adj_1582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19361_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__45932\,
            in1 => \N__50506\,
            in2 => \N__45926\,
            in3 => \N__50631\,
            lcout => n21968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19194_4_lut_3_lut_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55450\,
            in1 => \N__56505\,
            in2 => \_gnd_net_\,
            in3 => \N__56807\,
            lcout => \comm_spi.n14619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15244_2_lut_3_lut_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53951\,
            in1 => \N__45886\,
            in2 => \_gnd_net_\,
            in3 => \N__52365\,
            lcout => n14_adj_1578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19029_2_lut_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45854\,
            in2 => \_gnd_net_\,
            in3 => \N__56357\,
            lcout => n21270,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_238_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__46613\,
            in1 => \N__54824\,
            in2 => \N__49701\,
            in3 => \N__46586\,
            lcout => n12467,
            ltout => \n12467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46461\,
            in2 => \N__46550\,
            in3 => \N__46543\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_191_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__46523\,
            in1 => \N__46496\,
            in2 => \N__46465\,
            in3 => \N__46323\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21956_bdd_4_lut_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100100"
        )
    port map (
            in0 => \N__46880\,
            in1 => \N__46436\,
            in2 => \N__51873\,
            in3 => \N__49126\,
            lcout => n21959,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_102_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53950\,
            in1 => \N__46367\,
            in2 => \_gnd_net_\,
            in3 => \N__52364\,
            lcout => n14_adj_1577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46324\,
            in1 => \N__52174\,
            in2 => \_gnd_net_\,
            in3 => \N__47350\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__48418\,
            in1 => \N__49102\,
            in2 => \N__55700\,
            in3 => \N__46823\,
            lcout => OPEN,
            ltout => \n22208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22208_bdd_4_lut_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49103\,
            in1 => \N__46309\,
            in2 => \N__46292\,
            in3 => \N__46289\,
            lcout => OPEN,
            ltout => \n22211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1546664_i1_3_lut_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46262\,
            in2 => \N__47255\,
            in3 => \N__48676\,
            lcout => OPEN,
            ltout => \n30_adj_1518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54027\,
            in1 => \N__47246\,
            in2 => \N__47153\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57918\,
            ce => \N__47075\,
            sr => \N__46996\
        );

    \comm_cmd_1__bdd_4_lut_19375_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__46916\,
            in1 => \N__48414\,
            in2 => \N__46901\,
            in3 => \N__49101\,
            lcout => n21956,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_2_i26_3_lut_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46874\,
            in1 => \N__56362\,
            in2 => \_gnd_net_\,
            in3 => \N__46850\,
            lcout => n26_adj_1517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47376\,
            in1 => \N__46817\,
            in2 => \_gnd_net_\,
            in3 => \N__46690\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46796\,
            in1 => \N__47375\,
            in2 => \_gnd_net_\,
            in3 => \N__47506\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_188_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__46772\,
            in1 => \N__46745\,
            in2 => \N__46723\,
            in3 => \N__46689\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_5_i19_3_lut_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46670\,
            in1 => \N__46642\,
            in2 => \_gnd_net_\,
            in3 => \N__56338\,
            lcout => n19_adj_1497,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47377\,
            in1 => \N__47842\,
            in2 => \_gnd_net_\,
            in3 => \N__47701\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_134_Mux_7_i23_3_lut_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__51233\,
            in1 => \N__56337\,
            in2 => \_gnd_net_\,
            in3 => \N__47794\,
            lcout => n23_adj_1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_185_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47752\,
            in1 => \N__47732\,
            in2 => \N__47284\,
            in3 => \N__47700\,
            lcout => n20_adj_1596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15258_2_lut_3_lut_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47656\,
            in1 => \N__54076\,
            in2 => \_gnd_net_\,
            in3 => \N__52366\,
            lcout => n14_adj_1546,
            ltout => \n14_adj_1546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47380\,
            in1 => \_gnd_net_\,
            in2 => \N__47594\,
            in3 => \N__49153\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47575\,
            in1 => \N__47378\,
            in2 => \_gnd_net_\,
            in3 => \N__47551\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_180_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47531\,
            in1 => \N__47502\,
            in2 => \N__47486\,
            in3 => \N__47427\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47428\,
            in1 => \N__47461\,
            in2 => \_gnd_net_\,
            in3 => \N__47381\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47379\,
            in1 => \N__47326\,
            in2 => \_gnd_net_\,
            in3 => \N__47283\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49834\,
            in1 => \N__49372\,
            in2 => \N__51187\,
            in3 => \N__49275\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_135_Mux_7_i26_3_lut_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49253\,
            in1 => \N__56371\,
            in2 => \_gnd_net_\,
            in3 => \N__49229\,
            lcout => OPEN,
            ltout => \n26_adj_1500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18196_4_lut_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__56372\,
            in1 => \N__49205\,
            in2 => \N__49193\,
            in3 => \N__48415\,
            lcout => OPEN,
            ltout => \n20810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19454_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__49133\,
            in1 => \N__48730\,
            in2 => \N__49190\,
            in3 => \N__49121\,
            lcout => n22058,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18195_3_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48410\,
            in1 => \N__49180\,
            in2 => \_gnd_net_\,
            in3 => \N__49152\,
            lcout => n20809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011110011010"
        )
    port map (
            in0 => \N__48416\,
            in1 => \N__56373\,
            in2 => \N__48728\,
            in3 => \N__49123\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57953\,
            ce => \N__51443\,
            sr => \N__50405\
        );

    \comm_length_i1_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011110011111011"
        )
    port map (
            in0 => \N__49122\,
            in1 => \N__48677\,
            in2 => \N__56378\,
            in3 => \N__48417\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57953\,
            ce => \N__51443\,
            sr => \N__50405\
        );

    \i1_4_lut_adj_244_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47887\,
            in1 => \N__54308\,
            in2 => \N__47876\,
            in3 => \N__50684\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55237\,
            lcout => \comm_spi.data_tx_7__N_769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12253_3_lut_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__51435\,
            in1 => \N__52367\,
            in2 => \_gnd_net_\,
            in3 => \N__54912\,
            lcout => n14671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50262\,
            in2 => \_gnd_net_\,
            in3 => \N__50359\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57966\,
            ce => \N__50381\,
            sr => \N__50186\
        );

    \SIG_DDS.dds_state_i0_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__50396\,
            in1 => \N__50358\,
            in2 => \N__50390\,
            in3 => \N__50098\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57974\,
            ce => \N__50380\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.SCLK_27_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001010110001"
        )
    port map (
            in0 => \N__50361\,
            in1 => \N__50250\,
            in2 => \N__50026\,
            in3 => \N__50131\,
            lcout => \DDS_SCK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15030_2_lut_2_lut_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50009\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49978\,
            lcout => \CONT_SD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15087_2_lut_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54655\,
            in2 => \_gnd_net_\,
            in3 => \N__53562\,
            lcout => n17485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_224_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__51741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52304\,
            lcout => n20608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i46_2_lut_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51745\,
            in2 => \_gnd_net_\,
            in3 => \N__53955\,
            lcout => n23_adj_1501,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000000000"
        )
    port map (
            in0 => \N__53956\,
            in1 => \N__52302\,
            in2 => \N__51762\,
            in3 => \N__51690\,
            lcout => OPEN,
            ltout => \n21_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19152_4_lut_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101111111111"
        )
    port map (
            in0 => \N__52303\,
            in1 => \N__50828\,
            in2 => \N__50822\,
            in3 => \N__50819\,
            lcout => n18_adj_1633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12212_12213_set_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53327\,
            in1 => \N__53300\,
            in2 => \_gnd_net_\,
            in3 => \N__53279\,
            lcout => \comm_spi.n14630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57062\,
            ce => 'H',
            sr => \N__52526\
        );

    \comm_spi.i12200_3_lut_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53295\,
            in1 => \N__53277\,
            in2 => \_gnd_net_\,
            in3 => \N__53324\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19204_4_lut_3_lut_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50801\,
            in2 => \N__50804\,
            in3 => \N__56777\,
            lcout => \comm_spi.n22667\,
            ltout => \comm_spi.n22667_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12214_3_lut_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50795\,
            in2 => \N__50786\,
            in3 => \N__53306\,
            lcout => comm_rx_buf_0,
            ltout => \comm_rx_buf_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__50701\,
            in1 => \N__54723\,
            in2 => \N__50705\,
            in3 => \N__51298\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_2__bdd_4_lut_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__50662\,
            in1 => \N__50567\,
            in2 => \N__50969\,
            in3 => \N__50548\,
            lcout => n22172,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i5_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__51299\,
            in1 => \N__51042\,
            in2 => \N__54837\,
            in3 => \N__50968\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57867\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19189_4_lut_3_lut_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__53325\,
            in1 => \N__58135\,
            in2 => \_gnd_net_\,
            in3 => \N__56776\,
            lcout => \comm_spi.n22670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_290_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__54708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52368\,
            lcout => n12235,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_130_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__53787\,
            in1 => \N__52369\,
            in2 => \_gnd_net_\,
            in3 => \N__54709\,
            lcout => n19904,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i469_2_lut_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__51747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51688\,
            lcout => n2369,
            ltout => \n2369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19055_4_lut_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__52370\,
            in1 => \N__53788\,
            in2 => \N__50957\,
            in3 => \N__51746\,
            lcout => OPEN,
            ltout => \n21130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19149_4_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__53554\,
            in1 => \N__51611\,
            in2 => \N__50954\,
            in3 => \N__54710\,
            lcout => n14_adj_1506,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15091_2_lut_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53786\,
            in2 => \_gnd_net_\,
            in3 => \N__53553\,
            lcout => n3,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50932\,
            in2 => \N__50858\,
            in3 => \N__50850\,
            lcout => n19655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18885_2_lut_3_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51840\,
            in1 => \N__51689\,
            in2 => \_gnd_net_\,
            in3 => \N__53804\,
            lcout => n21129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18127_2_lut_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53805\,
            in2 => \_gnd_net_\,
            in3 => \N__53505\,
            lcout => n20740,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_178_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52420\,
            in2 => \_gnd_net_\,
            in3 => \N__53506\,
            lcout => OPEN,
            ltout => \n11363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_229_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__53806\,
            in1 => \N__51552\,
            in2 => \N__51593\,
            in3 => \N__54717\,
            lcout => n11935,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_88_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__53346\,
            in1 => \N__51551\,
            in2 => \N__51481\,
            in3 => \N__51455\,
            lcout => n11876,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i7_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__51266\,
            in1 => \N__54718\,
            in2 => \N__51407\,
            in3 => \N__51311\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i7_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51254\,
            lcout => buf_control_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57902\,
            ce => \N__51224\,
            sr => \N__51208\
        );

    \i15260_2_lut_3_lut_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__51181\,
            in1 => \N__53964\,
            in2 => \_gnd_net_\,
            in3 => \N__52412\,
            lcout => n14_adj_1548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i20_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53012\,
            in1 => \N__53254\,
            in2 => \N__51076\,
            in3 => \N__52088\,
            lcout => cmd_rdadctmp_20_adj_1430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57919\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15259_2_lut_3_lut_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__52493\,
            in1 => \N__53963\,
            in2 => \_gnd_net_\,
            in3 => \N__52411\,
            lcout => n14_adj_1547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19184_4_lut_3_lut_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56809\,
            in1 => \N__58055\,
            in2 => \_gnd_net_\,
            in3 => \N__56425\,
            lcout => \comm_spi.n22664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56506\,
            in2 => \_gnd_net_\,
            in3 => \N__56808\,
            lcout => \comm_spi.data_tx_7__N_767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i8_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53002\,
            in1 => \N__53179\,
            in2 => \N__52121\,
            in3 => \N__52143\,
            lcout => buf_adcdata_iac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19199_4_lut_3_lut_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56816\,
            in1 => \N__55020\,
            in2 => \_gnd_net_\,
            in3 => \N__55068\,
            lcout => \comm_spi.n22685\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i17_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__53003\,
            in1 => \N__52626\,
            in2 => \N__52120\,
            in3 => \N__52086\,
            lcout => cmd_rdadctmp_17_adj_1433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i18_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__52085\,
            in1 => \N__51885\,
            in2 => \N__52633\,
            in3 => \N__53007\,
            lcout => cmd_rdadctmp_18_adj_1432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i19_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__53004\,
            in1 => \N__53250\,
            in2 => \N__51890\,
            in3 => \N__52087\,
            lcout => cmd_rdadctmp_19_adj_1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i10_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53177\,
            in1 => \N__53005\,
            in2 => \N__51874\,
            in3 => \N__51889\,
            lcout => buf_adcdata_iac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19219_4_lut_3_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__58224\,
            in1 => \N__55272\,
            in2 => \_gnd_net_\,
            in3 => \N__56817\,
            lcout => \comm_spi.n22676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i11_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53178\,
            in1 => \N__53006\,
            in2 => \N__53255\,
            in3 => \N__53229\,
            lcout => buf_adcdata_iac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i9_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53176\,
            in1 => \N__53011\,
            in2 => \N__52634\,
            in3 => \N__52602\,
            lcout => buf_adcdata_iac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18953_2_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52583\,
            in2 => \_gnd_net_\,
            in3 => \N__56317\,
            lcout => n21230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__55027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56775\,
            lcout => \comm_spi.data_tx_7__N_793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19021_2_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__56313\,
            in1 => \N__52553\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n21297,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55127\,
            lcout => \comm_spi.DOUT_7__N_747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19209_4_lut_3_lut_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55386\,
            in1 => \N__55160\,
            in2 => \_gnd_net_\,
            in3 => \N__56745\,
            lcout => \comm_spi.n22682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__55318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56743\,
            lcout => \comm_spi.data_tx_7__N_787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56744\,
            lcout => \comm_spi.data_tx_7__N_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__56742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55510\,
            lcout => \comm_spi.data_tx_7__N_778\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_clear_311_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__54170\,
            in1 => \N__54913\,
            in2 => \_gnd_net_\,
            in3 => \N__53582\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57967\,
            ce => \N__54431\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_12228_12229_set_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__55187\,
            in1 => \N__55220\,
            in2 => \_gnd_net_\,
            in3 => \N__55201\,
            lcout => \comm_spi.n14646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57049\,
            ce => 'H',
            sr => \N__54416\
        );

    \mux_143_Mux_6_i4_3_lut_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__54407\,
            in1 => \N__54395\,
            in2 => \_gnd_net_\,
            in3 => \N__54368\,
            lcout => n4_adj_1585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6849_2_lut_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54028\,
            in2 => \_gnd_net_\,
            in3 => \N__53548\,
            lcout => n9270,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12212_12213_reset_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53326\,
            in1 => \N__53296\,
            in2 => \_gnd_net_\,
            in3 => \N__53278\,
            lcout => \comm_spi.n14631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57058\,
            ce => 'H',
            sr => \N__55106\
        );

    \comm_spi.imosi_44_12198_12199_set_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__58152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57891\,
            ce => 'H',
            sr => \N__55094\
        );

    \comm_spi.imosi_44_12198_12199_reset_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58153\,
            lcout => \comm_spi.n14617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57903\,
            ce => 'H',
            sr => \N__58097\
        );

    \comm_spi.imiso_83_12208_12209_set_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__56563\,
            in1 => \N__55412\,
            in2 => \_gnd_net_\,
            in3 => \N__55465\,
            lcout => \comm_spi.n14626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12208_12209_setC_net\,
            ce => 'H',
            sr => \N__56549\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55152\,
            in2 => \_gnd_net_\,
            in3 => \N__56836\,
            lcout => \comm_spi.data_tx_7__N_790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__55153\,
            in1 => \_gnd_net_\,
            in2 => \N__56853\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__56837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55123\,
            lcout => \comm_spi.DOUT_7__N_748\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58154\,
            in2 => \_gnd_net_\,
            in3 => \N__56835\,
            lcout => \comm_spi.imosi_N_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_12220_12221_reset_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55070\,
            in1 => \N__55043\,
            in2 => \_gnd_net_\,
            in3 => \N__56459\,
            lcout => \comm_spi.n14639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57012\,
            ce => 'H',
            sr => \N__55082\
        );

    \comm_spi.data_tx_i2_12220_12221_set_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55069\,
            in1 => \N__55039\,
            in2 => \_gnd_net_\,
            in3 => \N__56455\,
            lcout => \comm_spi.n14638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57017\,
            ce => 'H',
            sr => \N__55052\
        );

    \comm_spi.data_tx_i1_12216_12217_set_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56396\,
            in1 => \N__58085\,
            in2 => \_gnd_net_\,
            in3 => \N__57080\,
            lcout => \comm_spi.n14634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56917\,
            ce => 'H',
            sr => \N__54992\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56841\,
            lcout => \comm_spi.data_tx_7__N_773\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12194_12195_set_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58041\,
            lcout => \comm_spi.n14612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57961\,
            ce => 'H',
            sr => \N__56408\
        );

    \comm_spi.data_tx_i3_12224_12225_reset_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55393\,
            in1 => \N__55366\,
            in2 => \_gnd_net_\,
            in3 => \N__55339\,
            lcout => \comm_spi.n14643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56918\,
            ce => 'H',
            sr => \N__55325\
        );

    \comm_spi.i19214_4_lut_3_lut_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55218\,
            in1 => \N__55319\,
            in2 => \_gnd_net_\,
            in3 => \N__56749\,
            lcout => \comm_spi.n22679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55280\,
            in2 => \_gnd_net_\,
            in3 => \N__56747\,
            lcout => \comm_spi.data_tx_7__N_784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55511\,
            in2 => \_gnd_net_\,
            in3 => \N__56748\,
            lcout => \comm_spi.data_tx_7__N_768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__56746\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55246\,
            lcout => \comm_spi.data_tx_7__N_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19224_4_lut_3_lut_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55247\,
            in1 => \N__55653\,
            in2 => \_gnd_net_\,
            in3 => \N__56750\,
            lcout => \comm_spi.n22673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_12228_12229_reset_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55219\,
            in1 => \N__55202\,
            in2 => \_gnd_net_\,
            in3 => \N__55186\,
            lcout => \comm_spi.n14647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56997\,
            ce => 'H',
            sr => \N__55172\
        );

    \comm_spi.data_tx_i5_12232_12233_reset_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58237\,
            in1 => \N__58207\,
            in2 => \_gnd_net_\,
            in3 => \N__58192\,
            lcout => \comm_spi.n14651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57016\,
            ce => 'H',
            sr => \N__55604\
        );

    \i18943_2_lut_LC_20_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55592\,
            in2 => \_gnd_net_\,
            in3 => \N__56377\,
            lcout => n21204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12204_3_lut_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55478\,
            in1 => \N__55544\,
            in2 => \_gnd_net_\,
            in3 => \N__55520\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_12202_12203_reset_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__55538\,
            in1 => \N__55427\,
            in2 => \_gnd_net_\,
            in3 => \N__55477\,
            lcout => \comm_spi.n14621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12202_12203_resetC_net\,
            ce => 'H',
            sr => \N__56487\
        );

    \comm_spi.MISO_48_12202_12203_set_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55423\,
            in1 => \N__55534\,
            in2 => \_gnd_net_\,
            in3 => \N__55469\,
            lcout => \comm_spi.n14620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12202_12203_setC_net\,
            ce => 'H',
            sr => \N__56535\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56844\,
            lcout => \comm_spi.iclk_N_764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19229_4_lut_3_lut_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__56577\,
            in1 => \N__55497\,
            in2 => \_gnd_net_\,
            in3 => \N__56845\,
            lcout => \comm_spi.n22661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_12208_12209_reset_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__56564\,
            in1 => \N__55411\,
            in2 => \_gnd_net_\,
            in3 => \N__55476\,
            lcout => \comm_spi.n14627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12208_12209_resetC_net\,
            ce => 'H',
            sr => \N__56488\
        );

    \comm_spi.data_tx_i7_12205_12206_reset_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56584\,
            in1 => \N__55619\,
            in2 => \_gnd_net_\,
            in3 => \N__55685\,
            lcout => \comm_spi.n14624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56983\,
            ce => 'H',
            sr => \N__56489\
        );

    \comm_spi.data_tx_i7_12205_12206_set_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56585\,
            in1 => \N__55618\,
            in2 => \_gnd_net_\,
            in3 => \N__55684\,
            lcout => \comm_spi.n14623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56991\,
            ce => 'H',
            sr => \N__56542\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56513\,
            in2 => \_gnd_net_\,
            in3 => \N__56810\,
            lcout => \comm_spi.data_tx_7__N_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_12216_12217_reset_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56395\,
            in1 => \N__58084\,
            in2 => \_gnd_net_\,
            in3 => \N__57079\,
            lcout => \comm_spi.n14635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56910\,
            ce => 'H',
            sr => \N__56444\
        );

    \comm_spi.i12196_3_lut_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__57995\,
            in1 => \N__56432\,
            in2 => \_gnd_net_\,
            in3 => \N__56414\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58031\,
            in2 => \_gnd_net_\,
            in3 => \N__56832\,
            lcout => \comm_spi.iclk_N_763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19234_4_lut_3_lut_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__56632\,
            in1 => \N__56394\,
            in2 => \_gnd_net_\,
            in3 => \N__56833\,
            lcout => \comm_spi.n22688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19080_2_lut_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__56367\,
            in1 => \N__55712\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n21320,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12236_12237_reset_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55655\,
            in1 => \N__58181\,
            in2 => \_gnd_net_\,
            in3 => \N__55637\,
            lcout => \comm_spi.n14655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56911\,
            ce => 'H',
            sr => \N__55670\
        );

    \comm_spi.data_tx_i6_12236_12237_set_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55654\,
            in1 => \N__58177\,
            in2 => \_gnd_net_\,
            in3 => \N__55636\,
            lcout => \comm_spi.n14654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56987\,
            ce => 'H',
            sr => \N__58247\
        );

    \comm_spi.data_tx_i5_12232_12233_set_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58241\,
            in1 => \N__58208\,
            in2 => \_gnd_net_\,
            in3 => \N__58193\,
            lcout => \comm_spi.n14650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56996\,
            ce => 'H',
            sr => \N__58166\
        );

    \CONSTANT_ONE_LUT4_LC_22_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__58128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56842\,
            lcout => \comm_spi.imosi_N_754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56628\,
            in2 => \_gnd_net_\,
            in3 => \N__56843\,
            lcout => \comm_spi.data_tx_7__N_774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12190_12191_set_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__57186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57051\,
            ce => 'H',
            sr => \N__58067\
        );

    \comm_spi.iclk_40_12194_12195_reset_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__58054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57970\,
            ce => 'H',
            sr => \N__57440\
        );

    \comm_spi.data_tx_i0_12190_12191_reset_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__57237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__57040\,
            ce => 'H',
            sr => \N__56597\
        );

    \comm_spi.RESET_I_0_2_lut_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__56834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56633\,
            lcout => \comm_spi.data_tx_7__N_796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
