// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 28 2024 10:36:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "vdc_gen_clk" view "INTERFACE"

module vdc_gen_clk (
    DIVIDE,
    ICLK,
    OCLK);

    input [15:0] DIVIDE;
    input ICLK;
    output OCLK;

    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4236;
    wire N__4235;
    wire N__4234;
    wire N__4227;
    wire N__4226;
    wire N__4225;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4200;
    wire N__4199;
    wire N__4198;
    wire N__4191;
    wire N__4190;
    wire N__4189;
    wire N__4182;
    wire N__4181;
    wire N__4180;
    wire N__4173;
    wire N__4172;
    wire N__4171;
    wire N__4164;
    wire N__4163;
    wire N__4162;
    wire N__4155;
    wire N__4154;
    wire N__4153;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4137;
    wire N__4136;
    wire N__4135;
    wire N__4128;
    wire N__4127;
    wire N__4126;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4110;
    wire N__4109;
    wire N__4108;
    wire N__4101;
    wire N__4100;
    wire N__4099;
    wire N__4092;
    wire N__4091;
    wire N__4090;
    wire N__4073;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4055;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4043;
    wire N__4040;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4018;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4004;
    wire N__4001;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3986;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3932;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3922;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3823;
    wire N__3822;
    wire N__3821;
    wire N__3820;
    wire N__3819;
    wire N__3818;
    wire N__3817;
    wire N__3816;
    wire N__3815;
    wire N__3814;
    wire N__3813;
    wire N__3812;
    wire N__3811;
    wire N__3798;
    wire N__3795;
    wire N__3782;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3763;
    wire N__3762;
    wire N__3759;
    wire N__3758;
    wire N__3757;
    wire N__3756;
    wire N__3755;
    wire N__3754;
    wire N__3751;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3727;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3692;
    wire N__3691;
    wire N__3690;
    wire N__3689;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3681;
    wire N__3680;
    wire N__3679;
    wire N__3678;
    wire N__3677;
    wire N__3676;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3631;
    wire N__3626;
    wire N__3623;
    wire N__3618;
    wire N__3615;
    wire N__3614;
    wire N__3611;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3589;
    wire N__3586;
    wire N__3581;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3545;
    wire N__3542;
    wire N__3541;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3533;
    wire N__3530;
    wire N__3529;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3510;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3412;
    wire N__3411;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3403;
    wire N__3402;
    wire N__3399;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3372;
    wire N__3369;
    wire N__3364;
    wire N__3359;
    wire N__3356;
    wire N__3351;
    wire N__3344;
    wire N__3343;
    wire N__3342;
    wire N__3341;
    wire N__3340;
    wire N__3339;
    wire N__3338;
    wire N__3337;
    wire N__3336;
    wire N__3335;
    wire N__3334;
    wire N__3333;
    wire N__3330;
    wire N__3325;
    wire N__3324;
    wire N__3313;
    wire N__3304;
    wire N__3299;
    wire N__3298;
    wire N__3297;
    wire N__3294;
    wire N__3293;
    wire N__3288;
    wire N__3285;
    wire N__3278;
    wire N__3277;
    wire N__3276;
    wire N__3273;
    wire N__3272;
    wire N__3271;
    wire N__3268;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3250;
    wire N__3239;
    wire N__3236;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3221;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3206;
    wire N__3203;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3188;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3173;
    wire N__3170;
    wire N__3169;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3008;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2945;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2917;
    wire N__2912;
    wire N__2909;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2809;
    wire N__2808;
    wire N__2807;
    wire N__2806;
    wire N__2805;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2784;
    wire N__2783;
    wire N__2782;
    wire N__2781;
    wire N__2780;
    wire N__2779;
    wire N__2778;
    wire N__2777;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2773;
    wire N__2772;
    wire N__2771;
    wire N__2770;
    wire N__2769;
    wire N__2768;
    wire N__2761;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2728;
    wire N__2725;
    wire N__2724;
    wire N__2721;
    wire N__2720;
    wire N__2717;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2689;
    wire N__2682;
    wire N__2673;
    wire N__2656;
    wire N__2647;
    wire N__2640;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2608;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2549;
    wire N__2548;
    wire N__2545;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2535;
    wire N__2532;
    wire N__2527;
    wire N__2524;
    wire N__2521;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2506;
    wire N__2503;
    wire N__2500;
    wire N__2495;
    wire N__2492;
    wire N__2491;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2476;
    wire N__2473;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2458;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2435;
    wire N__2434;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2421;
    wire N__2416;
    wire N__2413;
    wire N__2410;
    wire N__2407;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2386;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2372;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2362;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2296;
    wire N__2293;
    wire N__2290;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2245;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2230;
    wire N__2227;
    wire N__2224;
    wire N__2221;
    wire N__2218;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2203;
    wire N__2200;
    wire N__2197;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2179;
    wire N__2176;
    wire N__2173;
    wire N__2168;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2143;
    wire N__2140;
    wire N__2137;
    wire N__2136;
    wire N__2133;
    wire N__2130;
    wire N__2127;
    wire N__2122;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2096;
    wire N__2093;
    wire N__2090;
    wire N__2089;
    wire N__2086;
    wire N__2083;
    wire N__2082;
    wire N__2079;
    wire N__2076;
    wire N__2073;
    wire N__2070;
    wire N__2065;
    wire N__2060;
    wire N__2057;
    wire N__2056;
    wire N__2053;
    wire N__2050;
    wire N__2049;
    wire N__2046;
    wire N__2043;
    wire N__2040;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2026;
    wire N__2023;
    wire N__2020;
    wire N__2015;
    wire N__2012;
    wire N__2009;
    wire N__2006;
    wire N__2005;
    wire N__2002;
    wire N__1999;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1981;
    wire N__1978;
    wire N__1975;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1946;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1931;
    wire N__1928;
    wire N__1927;
    wire N__1926;
    wire N__1923;
    wire N__1920;
    wire N__1917;
    wire N__1910;
    wire N__1907;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1877;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1865;
    wire N__1862;
    wire N__1859;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1851;
    wire N__1846;
    wire N__1843;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1798;
    wire N__1797;
    wire N__1794;
    wire N__1791;
    wire N__1788;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1769;
    wire N__1766;
    wire N__1763;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1751;
    wire N__1750;
    wire N__1747;
    wire N__1744;
    wire N__1739;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1699;
    wire N__1698;
    wire N__1695;
    wire N__1692;
    wire N__1689;
    wire N__1686;
    wire N__1681;
    wire N__1678;
    wire N__1675;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1625;
    wire N__1622;
    wire N__1619;
    wire VCCG0;
    wire GNDG0;
    wire DIVIDE_0_;
    wire bfn_1_9_0_;
    wire n16;
    wire n418;
    wire n15;
    wire n419;
    wire n14;
    wire n420;
    wire n13;
    wire DIVIDE_4_;
    wire n421;
    wire DIVIDE_5_;
    wire n422;
    wire n11;
    wire n423;
    wire n424;
    wire n425;
    wire n9;
    wire bfn_1_10_0_;
    wire DIVIDE_9_;
    wire n426;
    wire n427;
    wire n428;
    wire n5;
    wire n429;
    wire n4;
    wire n430;
    wire DIVIDE_14_;
    wire n431;
    wire n432;
    wire n7;
    wire OCLK;
    wire n10;
    wire DIVIDE_6_;
    wire n12;
    wire n3;
    wire DIVIDE_1_;
    wire n17;
    wire DIVIDE_7_;
    wire DIVIDE_2_;
    wire t0on_0;
    wire t0on_15_N_35_0;
    wire bfn_2_7_0_;
    wire t0on_1;
    wire t0on_15_N_35_1;
    wire n403;
    wire n404;
    wire t0on_3;
    wire t0on_15_N_35_3;
    wire n405;
    wire t0on_4;
    wire t0on_15_N_35_4;
    wire n406;
    wire t0on_5;
    wire t0on_15_N_35_5;
    wire n407;
    wire t0on_6;
    wire t0on_15_N_35_6;
    wire n408;
    wire n409;
    wire n410;
    wire t0on_8;
    wire t0on_15_N_35_8;
    wire bfn_2_8_0_;
    wire n411;
    wire n412;
    wire n413;
    wire n414;
    wire t0on_13;
    wire t0on_15_N_35_13;
    wire n415;
    wire n416;
    wire n417;
    wire bfn_2_9_0_;
    wire n388;
    wire n389;
    wire n390;
    wire n391;
    wire n392;
    wire n393;
    wire n394;
    wire n395;
    wire bfn_2_10_0_;
    wire n396;
    wire n397;
    wire n398;
    wire n399;
    wire n400;
    wire n401;
    wire CONSTANT_ONE_NET;
    wire n402;
    wire t0off_15_N_51_15;
    wire DIVIDE_11_;
    wire t0on_15_N_35_10;
    wire t0on_10;
    wire DIVIDE_3_;
    wire t0on_15_N_35_2;
    wire t0on_2;
    wire DIVIDE_13_;
    wire t0on_15_N_35_12;
    wire t0on_12;
    wire DIVIDE_8_;
    wire t0on_15_N_35_7;
    wire t0on_7;
    wire t0on_15;
    wire t0on_15_N_35_11;
    wire t0on_11;
    wire t0on_15_N_35_9;
    wire t0on_9;
    wire DIVIDE_15_;
    wire t0on_15_N_35_14;
    wire t0on_14;
    wire DIVIDE_12_;
    wire n6;
    wire DIVIDE_10_;
    wire n8;
    wire t0off_15_N_67_3;
    wire t0off_15_N_51_3;
    wire t0off_15_N_67_8;
    wire t0off_15_N_51_8;
    wire t0off_15_N_67_2;
    wire t0off_15_N_51_2;
    wire t0off_15_N_67_10;
    wire t0off_15_N_51_10;
    wire t0off_15_N_67_13;
    wire t0off_15_N_51_13;
    wire t0off_15_N_67_7;
    wire t0off_15_N_51_7;
    wire t0off_15_N_67_12;
    wire t0off_15_N_51_12;
    wire t0off_15_N_51_9;
    wire t0off_15_N_67_9;
    wire t0off_15_N_67_14;
    wire t0off_15_N_51_14;
    wire t0off_15_N_67_4;
    wire t0off_15_N_51_4;
    wire t0off_15_N_67_1;
    wire t0off_15_N_51_1;
    wire t0off_15_N_67_0;
    wire t0off_15_N_51_0;
    wire n26_adj_2;
    wire n27_adj_18;
    wire n28_adj_1;
    wire n447;
    wire n441_cascade_;
    wire n6_adj_3;
    wire n441;
    wire n386;
    wire div_state_1__N_88;
    wire div_state_0;
    wire t0off_12;
    wire t0off_2;
    wire t0off_7;
    wire t0off_10;
    wire n27_cascade_;
    wire n442;
    wire t0off_13;
    wire t0off_3;
    wire t0off_8;
    wire n26;
    wire t0off_14;
    wire t0off_15;
    wire t0off_9;
    wire n28;
    wire t0off_1;
    wire t0off_4;
    wire t0off_0;
    wire n444;
    wire t0off_15_N_67_5;
    wire t0off_15_N_51_5;
    wire t0off_5;
    wire t0off_15_N_67_6;
    wire t0off_15_N_51_6;
    wire t0off_6;
    wire t0off_15_N_67_11;
    wire div_state_1;
    wire t0off_15_N_51_11;
    wire t0off_11;
    wire ICLK;
    wire n307;
    wire _gnd_net_;

    IO_PAD ipInertedIOPad_DIVIDE_c_2_iopad (
            .OE(N__4245),
            .DIN(N__4244),
            .DOUT(N__4243),
            .PACKAGEPIN(DIVIDE[2]));
    defparam ipInertedIOPad_DIVIDE_c_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_2_preio (
            .PADOEN(N__4245),
            .PADOUT(N__4244),
            .PADIN(N__4243),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_2_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_10_iopad (
            .OE(N__4236),
            .DIN(N__4235),
            .DOUT(N__4234),
            .PACKAGEPIN(DIVIDE[10]));
    defparam ipInertedIOPad_DIVIDE_c_10_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_10_preio (
            .PADOEN(N__4236),
            .PADOUT(N__4235),
            .PADIN(N__4234),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_10_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_9_iopad (
            .OE(N__4227),
            .DIN(N__4226),
            .DOUT(N__4225),
            .PACKAGEPIN(DIVIDE[9]));
    defparam ipInertedIOPad_DIVIDE_c_9_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_9_preio (
            .PADOEN(N__4227),
            .PADOUT(N__4226),
            .PADIN(N__4225),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_9_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_5_iopad (
            .OE(N__4218),
            .DIN(N__4217),
            .DOUT(N__4216),
            .PACKAGEPIN(DIVIDE[5]));
    defparam ipInertedIOPad_DIVIDE_c_5_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_5_preio (
            .PADOEN(N__4218),
            .PADOUT(N__4217),
            .PADIN(N__4216),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_5_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_15_iopad (
            .OE(N__4209),
            .DIN(N__4208),
            .DOUT(N__4207),
            .PACKAGEPIN(DIVIDE[15]));
    defparam ipInertedIOPad_DIVIDE_c_15_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_15_preio (
            .PADOEN(N__4209),
            .PADOUT(N__4208),
            .PADIN(N__4207),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_15_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_11_iopad (
            .OE(N__4200),
            .DIN(N__4199),
            .DOUT(N__4198),
            .PACKAGEPIN(DIVIDE[11]));
    defparam ipInertedIOPad_DIVIDE_c_11_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_11_preio (
            .PADOEN(N__4200),
            .PADOUT(N__4199),
            .PADIN(N__4198),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_11_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_1_iopad (
            .OE(N__4191),
            .DIN(N__4190),
            .DOUT(N__4189),
            .PACKAGEPIN(DIVIDE[1]));
    defparam ipInertedIOPad_DIVIDE_c_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_1_preio (
            .PADOEN(N__4191),
            .PADOUT(N__4190),
            .PADIN(N__4189),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_1_),
            .DIN1());
    IO_PAD ipInertedIOPad_ICLK_iopad (
            .OE(N__4182),
            .DIN(N__4181),
            .DOUT(N__4180),
            .PACKAGEPIN(ICLK));
    defparam ipInertedIOPad_ICLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICLK_preio (
            .PADOEN(N__4182),
            .PADOUT(N__4181),
            .PADIN(N__4180),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICLK),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_8_iopad (
            .OE(N__4173),
            .DIN(N__4172),
            .DOUT(N__4171),
            .PACKAGEPIN(DIVIDE[8]));
    defparam ipInertedIOPad_DIVIDE_c_8_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_8_preio (
            .PADOEN(N__4173),
            .PADOUT(N__4172),
            .PADIN(N__4171),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_8_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_4_iopad (
            .OE(N__4164),
            .DIN(N__4163),
            .DOUT(N__4162),
            .PACKAGEPIN(DIVIDE[4]));
    defparam ipInertedIOPad_DIVIDE_c_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_4_preio (
            .PADOEN(N__4164),
            .PADOUT(N__4163),
            .PADIN(N__4162),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_4_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_12_iopad (
            .OE(N__4155),
            .DIN(N__4154),
            .DOUT(N__4153),
            .PACKAGEPIN(DIVIDE[12]));
    defparam ipInertedIOPad_DIVIDE_c_12_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_12_preio (
            .PADOEN(N__4155),
            .PADOUT(N__4154),
            .PADIN(N__4153),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_12_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_0_iopad (
            .OE(N__4146),
            .DIN(N__4145),
            .DOUT(N__4144),
            .PACKAGEPIN(DIVIDE[0]));
    defparam ipInertedIOPad_DIVIDE_c_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_0_preio (
            .PADOEN(N__4146),
            .PADOUT(N__4145),
            .PADIN(N__4144),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_0_),
            .DIN1());
    IO_PAD ipInertedIOPad_OCLK_iopad (
            .OE(N__4137),
            .DIN(N__4136),
            .DOUT(N__4135),
            .PACKAGEPIN(OCLK));
    defparam ipInertedIOPad_OCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_OCLK_preio (
            .PADOEN(N__4137),
            .PADOUT(N__4136),
            .PADIN(N__4135),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__1880),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_7_iopad (
            .OE(N__4128),
            .DIN(N__4127),
            .DOUT(N__4126),
            .PACKAGEPIN(DIVIDE[7]));
    defparam ipInertedIOPad_DIVIDE_c_7_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_7_preio (
            .PADOEN(N__4128),
            .PADOUT(N__4127),
            .PADIN(N__4126),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_7_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_3_iopad (
            .OE(N__4119),
            .DIN(N__4118),
            .DOUT(N__4117),
            .PACKAGEPIN(DIVIDE[3]));
    defparam ipInertedIOPad_DIVIDE_c_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_3_preio (
            .PADOEN(N__4119),
            .PADOUT(N__4118),
            .PADIN(N__4117),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_3_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_13_iopad (
            .OE(N__4110),
            .DIN(N__4109),
            .DOUT(N__4108),
            .PACKAGEPIN(DIVIDE[13]));
    defparam ipInertedIOPad_DIVIDE_c_13_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_13_preio (
            .PADOEN(N__4110),
            .PADOUT(N__4109),
            .PADIN(N__4108),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_13_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_6_iopad (
            .OE(N__4101),
            .DIN(N__4100),
            .DOUT(N__4099),
            .PACKAGEPIN(DIVIDE[6]));
    defparam ipInertedIOPad_DIVIDE_c_6_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_6_preio (
            .PADOEN(N__4101),
            .PADOUT(N__4100),
            .PADIN(N__4099),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_6_),
            .DIN1());
    IO_PAD ipInertedIOPad_DIVIDE_c_14_iopad (
            .OE(N__4092),
            .DIN(N__4091),
            .DOUT(N__4090),
            .PACKAGEPIN(DIVIDE[14]));
    defparam ipInertedIOPad_DIVIDE_c_14_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_DIVIDE_c_14_preio (
            .PADOEN(N__4092),
            .PADOUT(N__4091),
            .PADIN(N__4090),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(DIVIDE_14_),
            .DIN1());
    CascadeMux I__956 (
            .O(N__4073),
            .I(N__4069));
    InMux I__955 (
            .O(N__4072),
            .I(N__4066));
    InMux I__954 (
            .O(N__4069),
            .I(N__4063));
    LocalMux I__953 (
            .O(N__4066),
            .I(N__4060));
    LocalMux I__952 (
            .O(N__4063),
            .I(t0off_13));
    Odrv4 I__951 (
            .O(N__4060),
            .I(t0off_13));
    InMux I__950 (
            .O(N__4055),
            .I(N__4051));
    InMux I__949 (
            .O(N__4054),
            .I(N__4048));
    LocalMux I__948 (
            .O(N__4051),
            .I(N__4043));
    LocalMux I__947 (
            .O(N__4048),
            .I(N__4043));
    Odrv4 I__946 (
            .O(N__4043),
            .I(t0off_3));
    InMux I__945 (
            .O(N__4040),
            .I(N__4036));
    InMux I__944 (
            .O(N__4039),
            .I(N__4033));
    LocalMux I__943 (
            .O(N__4036),
            .I(N__4030));
    LocalMux I__942 (
            .O(N__4033),
            .I(t0off_8));
    Odrv4 I__941 (
            .O(N__4030),
            .I(t0off_8));
    InMux I__940 (
            .O(N__4025),
            .I(N__4022));
    LocalMux I__939 (
            .O(N__4022),
            .I(n26));
    InMux I__938 (
            .O(N__4019),
            .I(N__4015));
    InMux I__937 (
            .O(N__4018),
            .I(N__4012));
    LocalMux I__936 (
            .O(N__4015),
            .I(N__4009));
    LocalMux I__935 (
            .O(N__4012),
            .I(t0off_14));
    Odrv12 I__934 (
            .O(N__4009),
            .I(t0off_14));
    CascadeMux I__933 (
            .O(N__4004),
            .I(N__4001));
    InMux I__932 (
            .O(N__4001),
            .I(N__3997));
    InMux I__931 (
            .O(N__4000),
            .I(N__3994));
    LocalMux I__930 (
            .O(N__3997),
            .I(N__3991));
    LocalMux I__929 (
            .O(N__3994),
            .I(t0off_15));
    Odrv12 I__928 (
            .O(N__3991),
            .I(t0off_15));
    InMux I__927 (
            .O(N__3986),
            .I(N__3982));
    InMux I__926 (
            .O(N__3985),
            .I(N__3979));
    LocalMux I__925 (
            .O(N__3982),
            .I(N__3974));
    LocalMux I__924 (
            .O(N__3979),
            .I(N__3974));
    Odrv4 I__923 (
            .O(N__3974),
            .I(t0off_9));
    InMux I__922 (
            .O(N__3971),
            .I(N__3968));
    LocalMux I__921 (
            .O(N__3968),
            .I(n28));
    InMux I__920 (
            .O(N__3965),
            .I(N__3961));
    InMux I__919 (
            .O(N__3964),
            .I(N__3958));
    LocalMux I__918 (
            .O(N__3961),
            .I(N__3955));
    LocalMux I__917 (
            .O(N__3958),
            .I(t0off_1));
    Odrv4 I__916 (
            .O(N__3955),
            .I(t0off_1));
    CascadeMux I__915 (
            .O(N__3950),
            .I(N__3947));
    InMux I__914 (
            .O(N__3947),
            .I(N__3943));
    InMux I__913 (
            .O(N__3946),
            .I(N__3940));
    LocalMux I__912 (
            .O(N__3943),
            .I(N__3937));
    LocalMux I__911 (
            .O(N__3940),
            .I(t0off_4));
    Odrv4 I__910 (
            .O(N__3937),
            .I(t0off_4));
    InMux I__909 (
            .O(N__3932),
            .I(N__3928));
    InMux I__908 (
            .O(N__3931),
            .I(N__3925));
    LocalMux I__907 (
            .O(N__3928),
            .I(N__3922));
    LocalMux I__906 (
            .O(N__3925),
            .I(t0off_0));
    Odrv4 I__905 (
            .O(N__3922),
            .I(t0off_0));
    InMux I__904 (
            .O(N__3917),
            .I(N__3914));
    LocalMux I__903 (
            .O(N__3914),
            .I(n444));
    InMux I__902 (
            .O(N__3911),
            .I(N__3908));
    LocalMux I__901 (
            .O(N__3908),
            .I(N__3905));
    Odrv12 I__900 (
            .O(N__3905),
            .I(t0off_15_N_67_5));
    InMux I__899 (
            .O(N__3902),
            .I(N__3899));
    LocalMux I__898 (
            .O(N__3899),
            .I(N__3896));
    Span4Mux_h I__897 (
            .O(N__3896),
            .I(N__3893));
    Odrv4 I__896 (
            .O(N__3893),
            .I(t0off_15_N_51_5));
    InMux I__895 (
            .O(N__3890),
            .I(N__3886));
    CascadeMux I__894 (
            .O(N__3889),
            .I(N__3883));
    LocalMux I__893 (
            .O(N__3886),
            .I(N__3880));
    InMux I__892 (
            .O(N__3883),
            .I(N__3877));
    Span4Mux_h I__891 (
            .O(N__3880),
            .I(N__3872));
    LocalMux I__890 (
            .O(N__3877),
            .I(N__3872));
    Odrv4 I__889 (
            .O(N__3872),
            .I(t0off_5));
    InMux I__888 (
            .O(N__3869),
            .I(N__3866));
    LocalMux I__887 (
            .O(N__3866),
            .I(N__3863));
    Odrv12 I__886 (
            .O(N__3863),
            .I(t0off_15_N_67_6));
    InMux I__885 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__884 (
            .O(N__3857),
            .I(N__3854));
    Odrv12 I__883 (
            .O(N__3854),
            .I(t0off_15_N_51_6));
    InMux I__882 (
            .O(N__3851),
            .I(N__3848));
    LocalMux I__881 (
            .O(N__3848),
            .I(N__3844));
    InMux I__880 (
            .O(N__3847),
            .I(N__3841));
    Odrv12 I__879 (
            .O(N__3844),
            .I(t0off_6));
    LocalMux I__878 (
            .O(N__3841),
            .I(t0off_6));
    InMux I__877 (
            .O(N__3836),
            .I(N__3833));
    LocalMux I__876 (
            .O(N__3833),
            .I(N__3830));
    Span4Mux_h I__875 (
            .O(N__3830),
            .I(N__3827));
    Odrv4 I__874 (
            .O(N__3827),
            .I(t0off_15_N_67_11));
    InMux I__873 (
            .O(N__3824),
            .I(N__3798));
    InMux I__872 (
            .O(N__3823),
            .I(N__3798));
    InMux I__871 (
            .O(N__3822),
            .I(N__3798));
    InMux I__870 (
            .O(N__3821),
            .I(N__3798));
    InMux I__869 (
            .O(N__3820),
            .I(N__3798));
    InMux I__868 (
            .O(N__3819),
            .I(N__3798));
    InMux I__867 (
            .O(N__3818),
            .I(N__3795));
    InMux I__866 (
            .O(N__3817),
            .I(N__3782));
    InMux I__865 (
            .O(N__3816),
            .I(N__3782));
    InMux I__864 (
            .O(N__3815),
            .I(N__3782));
    InMux I__863 (
            .O(N__3814),
            .I(N__3782));
    InMux I__862 (
            .O(N__3813),
            .I(N__3782));
    InMux I__861 (
            .O(N__3812),
            .I(N__3782));
    InMux I__860 (
            .O(N__3811),
            .I(N__3777));
    LocalMux I__859 (
            .O(N__3798),
            .I(N__3774));
    LocalMux I__858 (
            .O(N__3795),
            .I(N__3771));
    LocalMux I__857 (
            .O(N__3782),
            .I(N__3768));
    InMux I__856 (
            .O(N__3781),
            .I(N__3763));
    InMux I__855 (
            .O(N__3780),
            .I(N__3763));
    LocalMux I__854 (
            .O(N__3777),
            .I(N__3759));
    Span4Mux_v I__853 (
            .O(N__3774),
            .I(N__3751));
    Span4Mux_v I__852 (
            .O(N__3771),
            .I(N__3744));
    Span4Mux_h I__851 (
            .O(N__3768),
            .I(N__3744));
    LocalMux I__850 (
            .O(N__3763),
            .I(N__3744));
    InMux I__849 (
            .O(N__3762),
            .I(N__3741));
    Span12Mux_v I__848 (
            .O(N__3759),
            .I(N__3738));
    InMux I__847 (
            .O(N__3758),
            .I(N__3727));
    InMux I__846 (
            .O(N__3757),
            .I(N__3727));
    InMux I__845 (
            .O(N__3756),
            .I(N__3727));
    InMux I__844 (
            .O(N__3755),
            .I(N__3727));
    InMux I__843 (
            .O(N__3754),
            .I(N__3727));
    Odrv4 I__842 (
            .O(N__3751),
            .I(div_state_1));
    Odrv4 I__841 (
            .O(N__3744),
            .I(div_state_1));
    LocalMux I__840 (
            .O(N__3741),
            .I(div_state_1));
    Odrv12 I__839 (
            .O(N__3738),
            .I(div_state_1));
    LocalMux I__838 (
            .O(N__3727),
            .I(div_state_1));
    InMux I__837 (
            .O(N__3716),
            .I(N__3713));
    LocalMux I__836 (
            .O(N__3713),
            .I(N__3710));
    Odrv12 I__835 (
            .O(N__3710),
            .I(t0off_15_N_51_11));
    InMux I__834 (
            .O(N__3707),
            .I(N__3704));
    LocalMux I__833 (
            .O(N__3704),
            .I(N__3700));
    InMux I__832 (
            .O(N__3703),
            .I(N__3697));
    Odrv12 I__831 (
            .O(N__3700),
            .I(t0off_11));
    LocalMux I__830 (
            .O(N__3697),
            .I(t0off_11));
    ClkMux I__829 (
            .O(N__3692),
            .I(N__3685));
    ClkMux I__828 (
            .O(N__3691),
            .I(N__3682));
    ClkMux I__827 (
            .O(N__3690),
            .I(N__3672));
    ClkMux I__826 (
            .O(N__3689),
            .I(N__3669));
    ClkMux I__825 (
            .O(N__3688),
            .I(N__3666));
    LocalMux I__824 (
            .O(N__3685),
            .I(N__3661));
    LocalMux I__823 (
            .O(N__3682),
            .I(N__3661));
    ClkMux I__822 (
            .O(N__3681),
            .I(N__3658));
    ClkMux I__821 (
            .O(N__3680),
            .I(N__3655));
    ClkMux I__820 (
            .O(N__3679),
            .I(N__3652));
    ClkMux I__819 (
            .O(N__3678),
            .I(N__3649));
    ClkMux I__818 (
            .O(N__3677),
            .I(N__3645));
    ClkMux I__817 (
            .O(N__3676),
            .I(N__3642));
    ClkMux I__816 (
            .O(N__3675),
            .I(N__3639));
    LocalMux I__815 (
            .O(N__3672),
            .I(N__3636));
    LocalMux I__814 (
            .O(N__3669),
            .I(N__3631));
    LocalMux I__813 (
            .O(N__3666),
            .I(N__3631));
    Span4Mux_h I__812 (
            .O(N__3661),
            .I(N__3626));
    LocalMux I__811 (
            .O(N__3658),
            .I(N__3626));
    LocalMux I__810 (
            .O(N__3655),
            .I(N__3623));
    LocalMux I__809 (
            .O(N__3652),
            .I(N__3618));
    LocalMux I__808 (
            .O(N__3649),
            .I(N__3618));
    ClkMux I__807 (
            .O(N__3648),
            .I(N__3615));
    LocalMux I__806 (
            .O(N__3645),
            .I(N__3611));
    LocalMux I__805 (
            .O(N__3642),
            .I(N__3606));
    LocalMux I__804 (
            .O(N__3639),
            .I(N__3606));
    Span4Mux_v I__803 (
            .O(N__3636),
            .I(N__3603));
    Span4Mux_v I__802 (
            .O(N__3631),
            .I(N__3600));
    Span4Mux_v I__801 (
            .O(N__3626),
            .I(N__3597));
    Span4Mux_v I__800 (
            .O(N__3623),
            .I(N__3594));
    Span4Mux_v I__799 (
            .O(N__3618),
            .I(N__3589));
    LocalMux I__798 (
            .O(N__3615),
            .I(N__3589));
    ClkMux I__797 (
            .O(N__3614),
            .I(N__3586));
    Span4Mux_v I__796 (
            .O(N__3611),
            .I(N__3581));
    Span4Mux_v I__795 (
            .O(N__3606),
            .I(N__3581));
    Span4Mux_h I__794 (
            .O(N__3603),
            .I(N__3568));
    Span4Mux_h I__793 (
            .O(N__3600),
            .I(N__3568));
    Span4Mux_v I__792 (
            .O(N__3597),
            .I(N__3568));
    Span4Mux_v I__791 (
            .O(N__3594),
            .I(N__3568));
    Span4Mux_v I__790 (
            .O(N__3589),
            .I(N__3568));
    LocalMux I__789 (
            .O(N__3586),
            .I(N__3568));
    Span4Mux_v I__788 (
            .O(N__3581),
            .I(N__3565));
    Span4Mux_h I__787 (
            .O(N__3568),
            .I(N__3562));
    Span4Mux_v I__786 (
            .O(N__3565),
            .I(N__3559));
    Span4Mux_v I__785 (
            .O(N__3562),
            .I(N__3556));
    Sp12to4 I__784 (
            .O(N__3559),
            .I(N__3553));
    Span4Mux_v I__783 (
            .O(N__3556),
            .I(N__3550));
    Odrv12 I__782 (
            .O(N__3553),
            .I(ICLK));
    Odrv4 I__781 (
            .O(N__3550),
            .I(ICLK));
    CEMux I__780 (
            .O(N__3545),
            .I(N__3542));
    LocalMux I__779 (
            .O(N__3542),
            .I(N__3537));
    CEMux I__778 (
            .O(N__3541),
            .I(N__3534));
    CEMux I__777 (
            .O(N__3540),
            .I(N__3530));
    Span4Mux_h I__776 (
            .O(N__3537),
            .I(N__3524));
    LocalMux I__775 (
            .O(N__3534),
            .I(N__3524));
    CEMux I__774 (
            .O(N__3533),
            .I(N__3521));
    LocalMux I__773 (
            .O(N__3530),
            .I(N__3518));
    CEMux I__772 (
            .O(N__3529),
            .I(N__3515));
    Span4Mux_h I__771 (
            .O(N__3524),
            .I(N__3510));
    LocalMux I__770 (
            .O(N__3521),
            .I(N__3510));
    Span4Mux_h I__769 (
            .O(N__3518),
            .I(N__3505));
    LocalMux I__768 (
            .O(N__3515),
            .I(N__3505));
    Span4Mux_h I__767 (
            .O(N__3510),
            .I(N__3502));
    Span4Mux_h I__766 (
            .O(N__3505),
            .I(N__3499));
    Odrv4 I__765 (
            .O(N__3502),
            .I(n307));
    Odrv4 I__764 (
            .O(N__3499),
            .I(n307));
    InMux I__763 (
            .O(N__3494),
            .I(N__3491));
    LocalMux I__762 (
            .O(N__3491),
            .I(N__3488));
    Span4Mux_h I__761 (
            .O(N__3488),
            .I(N__3485));
    Odrv4 I__760 (
            .O(N__3485),
            .I(n26_adj_2));
    InMux I__759 (
            .O(N__3482),
            .I(N__3479));
    LocalMux I__758 (
            .O(N__3479),
            .I(N__3476));
    Span4Mux_h I__757 (
            .O(N__3476),
            .I(N__3473));
    Odrv4 I__756 (
            .O(N__3473),
            .I(n27_adj_18));
    CascadeMux I__755 (
            .O(N__3470),
            .I(N__3467));
    InMux I__754 (
            .O(N__3467),
            .I(N__3464));
    LocalMux I__753 (
            .O(N__3464),
            .I(N__3461));
    Odrv4 I__752 (
            .O(N__3461),
            .I(n28_adj_1));
    InMux I__751 (
            .O(N__3458),
            .I(N__3455));
    LocalMux I__750 (
            .O(N__3455),
            .I(N__3452));
    Span4Mux_h I__749 (
            .O(N__3452),
            .I(N__3449));
    Odrv4 I__748 (
            .O(N__3449),
            .I(n447));
    CascadeMux I__747 (
            .O(N__3446),
            .I(n441_cascade_));
    CEMux I__746 (
            .O(N__3443),
            .I(N__3440));
    LocalMux I__745 (
            .O(N__3440),
            .I(N__3437));
    Span4Mux_v I__744 (
            .O(N__3437),
            .I(N__3434));
    Odrv4 I__743 (
            .O(N__3434),
            .I(n6_adj_3));
    InMux I__742 (
            .O(N__3431),
            .I(N__3428));
    LocalMux I__741 (
            .O(N__3428),
            .I(n441));
    SRMux I__740 (
            .O(N__3425),
            .I(N__3422));
    LocalMux I__739 (
            .O(N__3422),
            .I(N__3419));
    Span4Mux_h I__738 (
            .O(N__3419),
            .I(N__3416));
    Odrv4 I__737 (
            .O(N__3416),
            .I(n386));
    CEMux I__736 (
            .O(N__3413),
            .I(N__3408));
    CEMux I__735 (
            .O(N__3412),
            .I(N__3403));
    CEMux I__734 (
            .O(N__3411),
            .I(N__3399));
    LocalMux I__733 (
            .O(N__3408),
            .I(N__3395));
    CEMux I__732 (
            .O(N__3407),
            .I(N__3392));
    CEMux I__731 (
            .O(N__3406),
            .I(N__3389));
    LocalMux I__730 (
            .O(N__3403),
            .I(N__3386));
    InMux I__729 (
            .O(N__3402),
            .I(N__3383));
    LocalMux I__728 (
            .O(N__3399),
            .I(N__3380));
    CEMux I__727 (
            .O(N__3398),
            .I(N__3377));
    Span4Mux_v I__726 (
            .O(N__3395),
            .I(N__3372));
    LocalMux I__725 (
            .O(N__3392),
            .I(N__3372));
    LocalMux I__724 (
            .O(N__3389),
            .I(N__3369));
    Span4Mux_v I__723 (
            .O(N__3386),
            .I(N__3364));
    LocalMux I__722 (
            .O(N__3383),
            .I(N__3364));
    Span4Mux_v I__721 (
            .O(N__3380),
            .I(N__3359));
    LocalMux I__720 (
            .O(N__3377),
            .I(N__3359));
    Span4Mux_h I__719 (
            .O(N__3372),
            .I(N__3356));
    Span4Mux_h I__718 (
            .O(N__3369),
            .I(N__3351));
    Span4Mux_h I__717 (
            .O(N__3364),
            .I(N__3351));
    Odrv4 I__716 (
            .O(N__3359),
            .I(div_state_1__N_88));
    Odrv4 I__715 (
            .O(N__3356),
            .I(div_state_1__N_88));
    Odrv4 I__714 (
            .O(N__3351),
            .I(div_state_1__N_88));
    InMux I__713 (
            .O(N__3344),
            .I(N__3330));
    InMux I__712 (
            .O(N__3343),
            .I(N__3325));
    InMux I__711 (
            .O(N__3342),
            .I(N__3325));
    InMux I__710 (
            .O(N__3341),
            .I(N__3313));
    InMux I__709 (
            .O(N__3340),
            .I(N__3313));
    InMux I__708 (
            .O(N__3339),
            .I(N__3313));
    InMux I__707 (
            .O(N__3338),
            .I(N__3313));
    InMux I__706 (
            .O(N__3337),
            .I(N__3313));
    InMux I__705 (
            .O(N__3336),
            .I(N__3304));
    InMux I__704 (
            .O(N__3335),
            .I(N__3304));
    InMux I__703 (
            .O(N__3334),
            .I(N__3304));
    InMux I__702 (
            .O(N__3333),
            .I(N__3304));
    LocalMux I__701 (
            .O(N__3330),
            .I(N__3299));
    LocalMux I__700 (
            .O(N__3325),
            .I(N__3299));
    CascadeMux I__699 (
            .O(N__3324),
            .I(N__3294));
    LocalMux I__698 (
            .O(N__3313),
            .I(N__3288));
    LocalMux I__697 (
            .O(N__3304),
            .I(N__3288));
    Span4Mux_v I__696 (
            .O(N__3299),
            .I(N__3285));
    InMux I__695 (
            .O(N__3298),
            .I(N__3278));
    InMux I__694 (
            .O(N__3297),
            .I(N__3278));
    InMux I__693 (
            .O(N__3294),
            .I(N__3278));
    CascadeMux I__692 (
            .O(N__3293),
            .I(N__3273));
    Span4Mux_h I__691 (
            .O(N__3288),
            .I(N__3268));
    Sp12to4 I__690 (
            .O(N__3285),
            .I(N__3263));
    LocalMux I__689 (
            .O(N__3278),
            .I(N__3263));
    InMux I__688 (
            .O(N__3277),
            .I(N__3260));
    InMux I__687 (
            .O(N__3276),
            .I(N__3257));
    InMux I__686 (
            .O(N__3273),
            .I(N__3250));
    InMux I__685 (
            .O(N__3272),
            .I(N__3250));
    InMux I__684 (
            .O(N__3271),
            .I(N__3250));
    Odrv4 I__683 (
            .O(N__3268),
            .I(div_state_0));
    Odrv12 I__682 (
            .O(N__3263),
            .I(div_state_0));
    LocalMux I__681 (
            .O(N__3260),
            .I(div_state_0));
    LocalMux I__680 (
            .O(N__3257),
            .I(div_state_0));
    LocalMux I__679 (
            .O(N__3250),
            .I(div_state_0));
    InMux I__678 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__677 (
            .O(N__3236),
            .I(N__3232));
    InMux I__676 (
            .O(N__3235),
            .I(N__3229));
    Span4Mux_v I__675 (
            .O(N__3232),
            .I(N__3226));
    LocalMux I__674 (
            .O(N__3229),
            .I(t0off_12));
    Odrv4 I__673 (
            .O(N__3226),
            .I(t0off_12));
    InMux I__672 (
            .O(N__3221),
            .I(N__3217));
    InMux I__671 (
            .O(N__3220),
            .I(N__3214));
    LocalMux I__670 (
            .O(N__3217),
            .I(N__3211));
    LocalMux I__669 (
            .O(N__3214),
            .I(t0off_2));
    Odrv4 I__668 (
            .O(N__3211),
            .I(t0off_2));
    CascadeMux I__667 (
            .O(N__3206),
            .I(N__3203));
    InMux I__666 (
            .O(N__3203),
            .I(N__3199));
    InMux I__665 (
            .O(N__3202),
            .I(N__3196));
    LocalMux I__664 (
            .O(N__3199),
            .I(N__3193));
    LocalMux I__663 (
            .O(N__3196),
            .I(t0off_7));
    Odrv4 I__662 (
            .O(N__3193),
            .I(t0off_7));
    InMux I__661 (
            .O(N__3188),
            .I(N__3184));
    InMux I__660 (
            .O(N__3187),
            .I(N__3181));
    LocalMux I__659 (
            .O(N__3184),
            .I(N__3178));
    LocalMux I__658 (
            .O(N__3181),
            .I(t0off_10));
    Odrv4 I__657 (
            .O(N__3178),
            .I(t0off_10));
    CascadeMux I__656 (
            .O(N__3173),
            .I(n27_cascade_));
    InMux I__655 (
            .O(N__3170),
            .I(N__3164));
    InMux I__654 (
            .O(N__3169),
            .I(N__3164));
    LocalMux I__653 (
            .O(N__3164),
            .I(n442));
    InMux I__652 (
            .O(N__3161),
            .I(N__3158));
    LocalMux I__651 (
            .O(N__3158),
            .I(N__3155));
    Span4Mux_h I__650 (
            .O(N__3155),
            .I(N__3152));
    Odrv4 I__649 (
            .O(N__3152),
            .I(t0off_15_N_67_13));
    InMux I__648 (
            .O(N__3149),
            .I(N__3146));
    LocalMux I__647 (
            .O(N__3146),
            .I(t0off_15_N_51_13));
    InMux I__646 (
            .O(N__3143),
            .I(N__3140));
    LocalMux I__645 (
            .O(N__3140),
            .I(N__3137));
    Odrv4 I__644 (
            .O(N__3137),
            .I(t0off_15_N_67_7));
    InMux I__643 (
            .O(N__3134),
            .I(N__3131));
    LocalMux I__642 (
            .O(N__3131),
            .I(t0off_15_N_51_7));
    InMux I__641 (
            .O(N__3128),
            .I(N__3125));
    LocalMux I__640 (
            .O(N__3125),
            .I(N__3122));
    Odrv12 I__639 (
            .O(N__3122),
            .I(t0off_15_N_67_12));
    InMux I__638 (
            .O(N__3119),
            .I(N__3116));
    LocalMux I__637 (
            .O(N__3116),
            .I(t0off_15_N_51_12));
    InMux I__636 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__635 (
            .O(N__3110),
            .I(t0off_15_N_51_9));
    InMux I__634 (
            .O(N__3107),
            .I(N__3104));
    LocalMux I__633 (
            .O(N__3104),
            .I(N__3101));
    Odrv4 I__632 (
            .O(N__3101),
            .I(t0off_15_N_67_9));
    InMux I__631 (
            .O(N__3098),
            .I(N__3095));
    LocalMux I__630 (
            .O(N__3095),
            .I(N__3092));
    Odrv12 I__629 (
            .O(N__3092),
            .I(t0off_15_N_67_14));
    InMux I__628 (
            .O(N__3089),
            .I(N__3086));
    LocalMux I__627 (
            .O(N__3086),
            .I(t0off_15_N_51_14));
    InMux I__626 (
            .O(N__3083),
            .I(N__3080));
    LocalMux I__625 (
            .O(N__3080),
            .I(N__3077));
    Span4Mux_v I__624 (
            .O(N__3077),
            .I(N__3074));
    Odrv4 I__623 (
            .O(N__3074),
            .I(t0off_15_N_67_4));
    InMux I__622 (
            .O(N__3071),
            .I(N__3068));
    LocalMux I__621 (
            .O(N__3068),
            .I(t0off_15_N_51_4));
    InMux I__620 (
            .O(N__3065),
            .I(N__3062));
    LocalMux I__619 (
            .O(N__3062),
            .I(N__3059));
    Span4Mux_v I__618 (
            .O(N__3059),
            .I(N__3056));
    Odrv4 I__617 (
            .O(N__3056),
            .I(t0off_15_N_67_1));
    InMux I__616 (
            .O(N__3053),
            .I(N__3050));
    LocalMux I__615 (
            .O(N__3050),
            .I(t0off_15_N_51_1));
    InMux I__614 (
            .O(N__3047),
            .I(N__3044));
    LocalMux I__613 (
            .O(N__3044),
            .I(N__3041));
    Span4Mux_h I__612 (
            .O(N__3041),
            .I(N__3038));
    Odrv4 I__611 (
            .O(N__3038),
            .I(t0off_15_N_67_0));
    InMux I__610 (
            .O(N__3035),
            .I(N__3032));
    LocalMux I__609 (
            .O(N__3032),
            .I(t0off_15_N_51_0));
    InMux I__608 (
            .O(N__3029),
            .I(N__3026));
    LocalMux I__607 (
            .O(N__3026),
            .I(t0on_15_N_35_9));
    CascadeMux I__606 (
            .O(N__3023),
            .I(N__3020));
    InMux I__605 (
            .O(N__3020),
            .I(N__3016));
    InMux I__604 (
            .O(N__3019),
            .I(N__3013));
    LocalMux I__603 (
            .O(N__3016),
            .I(t0on_9));
    LocalMux I__602 (
            .O(N__3013),
            .I(t0on_9));
    InMux I__601 (
            .O(N__3008),
            .I(N__3004));
    InMux I__600 (
            .O(N__3007),
            .I(N__3001));
    LocalMux I__599 (
            .O(N__3004),
            .I(N__2998));
    LocalMux I__598 (
            .O(N__3001),
            .I(N__2995));
    Span4Mux_v I__597 (
            .O(N__2998),
            .I(N__2991));
    Span4Mux_v I__596 (
            .O(N__2995),
            .I(N__2988));
    InMux I__595 (
            .O(N__2994),
            .I(N__2985));
    Sp12to4 I__594 (
            .O(N__2991),
            .I(N__2978));
    Sp12to4 I__593 (
            .O(N__2988),
            .I(N__2978));
    LocalMux I__592 (
            .O(N__2985),
            .I(N__2978));
    Odrv12 I__591 (
            .O(N__2978),
            .I(DIVIDE_15_));
    InMux I__590 (
            .O(N__2975),
            .I(N__2972));
    LocalMux I__589 (
            .O(N__2972),
            .I(t0on_15_N_35_14));
    InMux I__588 (
            .O(N__2969),
            .I(N__2965));
    InMux I__587 (
            .O(N__2968),
            .I(N__2962));
    LocalMux I__586 (
            .O(N__2965),
            .I(t0on_14));
    LocalMux I__585 (
            .O(N__2962),
            .I(t0on_14));
    InMux I__584 (
            .O(N__2957),
            .I(N__2953));
    InMux I__583 (
            .O(N__2956),
            .I(N__2950));
    LocalMux I__582 (
            .O(N__2953),
            .I(N__2945));
    LocalMux I__581 (
            .O(N__2950),
            .I(N__2945));
    Span4Mux_v I__580 (
            .O(N__2945),
            .I(N__2941));
    InMux I__579 (
            .O(N__2944),
            .I(N__2938));
    Sp12to4 I__578 (
            .O(N__2941),
            .I(N__2933));
    LocalMux I__577 (
            .O(N__2938),
            .I(N__2933));
    Odrv12 I__576 (
            .O(N__2933),
            .I(DIVIDE_12_));
    InMux I__575 (
            .O(N__2930),
            .I(N__2927));
    LocalMux I__574 (
            .O(N__2927),
            .I(N__2924));
    Span4Mux_v I__573 (
            .O(N__2924),
            .I(N__2921));
    Odrv4 I__572 (
            .O(N__2921),
            .I(n6));
    InMux I__571 (
            .O(N__2918),
            .I(N__2912));
    InMux I__570 (
            .O(N__2917),
            .I(N__2912));
    LocalMux I__569 (
            .O(N__2912),
            .I(N__2909));
    Span4Mux_v I__568 (
            .O(N__2909),
            .I(N__2905));
    InMux I__567 (
            .O(N__2908),
            .I(N__2902));
    Sp12to4 I__566 (
            .O(N__2905),
            .I(N__2897));
    LocalMux I__565 (
            .O(N__2902),
            .I(N__2897));
    Odrv12 I__564 (
            .O(N__2897),
            .I(DIVIDE_10_));
    CascadeMux I__563 (
            .O(N__2894),
            .I(N__2891));
    InMux I__562 (
            .O(N__2891),
            .I(N__2888));
    LocalMux I__561 (
            .O(N__2888),
            .I(N__2885));
    Span4Mux_v I__560 (
            .O(N__2885),
            .I(N__2882));
    Odrv4 I__559 (
            .O(N__2882),
            .I(n8));
    InMux I__558 (
            .O(N__2879),
            .I(N__2876));
    LocalMux I__557 (
            .O(N__2876),
            .I(N__2873));
    Odrv12 I__556 (
            .O(N__2873),
            .I(t0off_15_N_67_3));
    InMux I__555 (
            .O(N__2870),
            .I(N__2867));
    LocalMux I__554 (
            .O(N__2867),
            .I(t0off_15_N_51_3));
    InMux I__553 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__552 (
            .O(N__2861),
            .I(N__2858));
    Span4Mux_v I__551 (
            .O(N__2858),
            .I(N__2855));
    Odrv4 I__550 (
            .O(N__2855),
            .I(t0off_15_N_67_8));
    InMux I__549 (
            .O(N__2852),
            .I(N__2849));
    LocalMux I__548 (
            .O(N__2849),
            .I(t0off_15_N_51_8));
    InMux I__547 (
            .O(N__2846),
            .I(N__2843));
    LocalMux I__546 (
            .O(N__2843),
            .I(N__2840));
    Odrv4 I__545 (
            .O(N__2840),
            .I(t0off_15_N_67_2));
    InMux I__544 (
            .O(N__2837),
            .I(N__2834));
    LocalMux I__543 (
            .O(N__2834),
            .I(t0off_15_N_51_2));
    CascadeMux I__542 (
            .O(N__2831),
            .I(N__2828));
    InMux I__541 (
            .O(N__2828),
            .I(N__2825));
    LocalMux I__540 (
            .O(N__2825),
            .I(N__2822));
    Span4Mux_v I__539 (
            .O(N__2822),
            .I(N__2819));
    Odrv4 I__538 (
            .O(N__2819),
            .I(t0off_15_N_67_10));
    InMux I__537 (
            .O(N__2816),
            .I(N__2813));
    LocalMux I__536 (
            .O(N__2813),
            .I(t0off_15_N_51_10));
    CascadeMux I__535 (
            .O(N__2810),
            .I(N__2801));
    CascadeMux I__534 (
            .O(N__2809),
            .I(N__2798));
    CascadeMux I__533 (
            .O(N__2808),
            .I(N__2795));
    CascadeMux I__532 (
            .O(N__2807),
            .I(N__2791));
    CascadeMux I__531 (
            .O(N__2806),
            .I(N__2788));
    CascadeMux I__530 (
            .O(N__2805),
            .I(N__2785));
    InMux I__529 (
            .O(N__2804),
            .I(N__2761));
    InMux I__528 (
            .O(N__2801),
            .I(N__2761));
    InMux I__527 (
            .O(N__2798),
            .I(N__2761));
    InMux I__526 (
            .O(N__2795),
            .I(N__2750));
    InMux I__525 (
            .O(N__2794),
            .I(N__2750));
    InMux I__524 (
            .O(N__2791),
            .I(N__2750));
    InMux I__523 (
            .O(N__2788),
            .I(N__2750));
    InMux I__522 (
            .O(N__2785),
            .I(N__2750));
    CascadeMux I__521 (
            .O(N__2784),
            .I(N__2747));
    CascadeMux I__520 (
            .O(N__2783),
            .I(N__2744));
    CascadeMux I__519 (
            .O(N__2782),
            .I(N__2741));
    CascadeMux I__518 (
            .O(N__2781),
            .I(N__2738));
    CascadeMux I__517 (
            .O(N__2780),
            .I(N__2735));
    CascadeMux I__516 (
            .O(N__2779),
            .I(N__2732));
    CascadeMux I__515 (
            .O(N__2778),
            .I(N__2729));
    CascadeMux I__514 (
            .O(N__2777),
            .I(N__2725));
    CascadeMux I__513 (
            .O(N__2776),
            .I(N__2721));
    CascadeMux I__512 (
            .O(N__2775),
            .I(N__2717));
    CascadeMux I__511 (
            .O(N__2774),
            .I(N__2713));
    CascadeMux I__510 (
            .O(N__2773),
            .I(N__2710));
    CascadeMux I__509 (
            .O(N__2772),
            .I(N__2706));
    CascadeMux I__508 (
            .O(N__2771),
            .I(N__2703));
    CascadeMux I__507 (
            .O(N__2770),
            .I(N__2700));
    CascadeMux I__506 (
            .O(N__2769),
            .I(N__2697));
    CascadeMux I__505 (
            .O(N__2768),
            .I(N__2694));
    LocalMux I__504 (
            .O(N__2761),
            .I(N__2689));
    LocalMux I__503 (
            .O(N__2750),
            .I(N__2689));
    InMux I__502 (
            .O(N__2747),
            .I(N__2682));
    InMux I__501 (
            .O(N__2744),
            .I(N__2682));
    InMux I__500 (
            .O(N__2741),
            .I(N__2682));
    InMux I__499 (
            .O(N__2738),
            .I(N__2673));
    InMux I__498 (
            .O(N__2735),
            .I(N__2673));
    InMux I__497 (
            .O(N__2732),
            .I(N__2673));
    InMux I__496 (
            .O(N__2729),
            .I(N__2673));
    InMux I__495 (
            .O(N__2728),
            .I(N__2656));
    InMux I__494 (
            .O(N__2725),
            .I(N__2656));
    InMux I__493 (
            .O(N__2724),
            .I(N__2656));
    InMux I__492 (
            .O(N__2721),
            .I(N__2656));
    InMux I__491 (
            .O(N__2720),
            .I(N__2656));
    InMux I__490 (
            .O(N__2717),
            .I(N__2656));
    InMux I__489 (
            .O(N__2716),
            .I(N__2656));
    InMux I__488 (
            .O(N__2713),
            .I(N__2656));
    InMux I__487 (
            .O(N__2710),
            .I(N__2647));
    InMux I__486 (
            .O(N__2709),
            .I(N__2647));
    InMux I__485 (
            .O(N__2706),
            .I(N__2647));
    InMux I__484 (
            .O(N__2703),
            .I(N__2647));
    InMux I__483 (
            .O(N__2700),
            .I(N__2640));
    InMux I__482 (
            .O(N__2697),
            .I(N__2640));
    InMux I__481 (
            .O(N__2694),
            .I(N__2640));
    Span4Mux_v I__480 (
            .O(N__2689),
            .I(N__2627));
    LocalMux I__479 (
            .O(N__2682),
            .I(N__2627));
    LocalMux I__478 (
            .O(N__2673),
            .I(N__2627));
    LocalMux I__477 (
            .O(N__2656),
            .I(N__2627));
    LocalMux I__476 (
            .O(N__2647),
            .I(N__2627));
    LocalMux I__475 (
            .O(N__2640),
            .I(N__2627));
    Span4Mux_v I__474 (
            .O(N__2627),
            .I(N__2624));
    Odrv4 I__473 (
            .O(N__2624),
            .I(CONSTANT_ONE_NET));
    InMux I__472 (
            .O(N__2621),
            .I(n402));
    CascadeMux I__471 (
            .O(N__2618),
            .I(N__2615));
    InMux I__470 (
            .O(N__2615),
            .I(N__2612));
    LocalMux I__469 (
            .O(N__2612),
            .I(t0off_15_N_51_15));
    CascadeMux I__468 (
            .O(N__2609),
            .I(N__2604));
    InMux I__467 (
            .O(N__2608),
            .I(N__2601));
    InMux I__466 (
            .O(N__2607),
            .I(N__2598));
    InMux I__465 (
            .O(N__2604),
            .I(N__2595));
    LocalMux I__464 (
            .O(N__2601),
            .I(N__2592));
    LocalMux I__463 (
            .O(N__2598),
            .I(N__2587));
    LocalMux I__462 (
            .O(N__2595),
            .I(N__2587));
    Span4Mux_v I__461 (
            .O(N__2592),
            .I(N__2584));
    Sp12to4 I__460 (
            .O(N__2587),
            .I(N__2581));
    Span4Mux_h I__459 (
            .O(N__2584),
            .I(N__2578));
    Span12Mux_v I__458 (
            .O(N__2581),
            .I(N__2575));
    Span4Mux_v I__457 (
            .O(N__2578),
            .I(N__2572));
    Odrv12 I__456 (
            .O(N__2575),
            .I(DIVIDE_11_));
    Odrv4 I__455 (
            .O(N__2572),
            .I(DIVIDE_11_));
    InMux I__454 (
            .O(N__2567),
            .I(N__2564));
    LocalMux I__453 (
            .O(N__2564),
            .I(t0on_15_N_35_10));
    InMux I__452 (
            .O(N__2561),
            .I(N__2557));
    InMux I__451 (
            .O(N__2560),
            .I(N__2554));
    LocalMux I__450 (
            .O(N__2557),
            .I(t0on_10));
    LocalMux I__449 (
            .O(N__2554),
            .I(t0on_10));
    CascadeMux I__448 (
            .O(N__2549),
            .I(N__2545));
    InMux I__447 (
            .O(N__2548),
            .I(N__2541));
    InMux I__446 (
            .O(N__2545),
            .I(N__2538));
    InMux I__445 (
            .O(N__2544),
            .I(N__2535));
    LocalMux I__444 (
            .O(N__2541),
            .I(N__2532));
    LocalMux I__443 (
            .O(N__2538),
            .I(N__2527));
    LocalMux I__442 (
            .O(N__2535),
            .I(N__2527));
    Sp12to4 I__441 (
            .O(N__2532),
            .I(N__2524));
    Span4Mux_v I__440 (
            .O(N__2527),
            .I(N__2521));
    Span12Mux_v I__439 (
            .O(N__2524),
            .I(N__2516));
    Sp12to4 I__438 (
            .O(N__2521),
            .I(N__2516));
    Odrv12 I__437 (
            .O(N__2516),
            .I(DIVIDE_3_));
    InMux I__436 (
            .O(N__2513),
            .I(N__2510));
    LocalMux I__435 (
            .O(N__2510),
            .I(t0on_15_N_35_2));
    InMux I__434 (
            .O(N__2507),
            .I(N__2503));
    InMux I__433 (
            .O(N__2506),
            .I(N__2500));
    LocalMux I__432 (
            .O(N__2503),
            .I(t0on_2));
    LocalMux I__431 (
            .O(N__2500),
            .I(t0on_2));
    InMux I__430 (
            .O(N__2495),
            .I(N__2492));
    LocalMux I__429 (
            .O(N__2492),
            .I(N__2487));
    InMux I__428 (
            .O(N__2491),
            .I(N__2484));
    InMux I__427 (
            .O(N__2490),
            .I(N__2481));
    Span4Mux_v I__426 (
            .O(N__2487),
            .I(N__2476));
    LocalMux I__425 (
            .O(N__2484),
            .I(N__2476));
    LocalMux I__424 (
            .O(N__2481),
            .I(N__2473));
    Span4Mux_v I__423 (
            .O(N__2476),
            .I(N__2470));
    Sp12to4 I__422 (
            .O(N__2473),
            .I(N__2467));
    Span4Mux_h I__421 (
            .O(N__2470),
            .I(N__2464));
    Span12Mux_v I__420 (
            .O(N__2467),
            .I(N__2461));
    Span4Mux_v I__419 (
            .O(N__2464),
            .I(N__2458));
    Odrv12 I__418 (
            .O(N__2461),
            .I(DIVIDE_13_));
    Odrv4 I__417 (
            .O(N__2458),
            .I(DIVIDE_13_));
    InMux I__416 (
            .O(N__2453),
            .I(N__2450));
    LocalMux I__415 (
            .O(N__2450),
            .I(t0on_15_N_35_12));
    InMux I__414 (
            .O(N__2447),
            .I(N__2443));
    InMux I__413 (
            .O(N__2446),
            .I(N__2440));
    LocalMux I__412 (
            .O(N__2443),
            .I(t0on_12));
    LocalMux I__411 (
            .O(N__2440),
            .I(t0on_12));
    InMux I__410 (
            .O(N__2435),
            .I(N__2430));
    InMux I__409 (
            .O(N__2434),
            .I(N__2427));
    InMux I__408 (
            .O(N__2433),
            .I(N__2424));
    LocalMux I__407 (
            .O(N__2430),
            .I(N__2421));
    LocalMux I__406 (
            .O(N__2427),
            .I(N__2416));
    LocalMux I__405 (
            .O(N__2424),
            .I(N__2416));
    Span4Mux_v I__404 (
            .O(N__2421),
            .I(N__2413));
    Span4Mux_v I__403 (
            .O(N__2416),
            .I(N__2410));
    Sp12to4 I__402 (
            .O(N__2413),
            .I(N__2407));
    Span4Mux_v I__401 (
            .O(N__2410),
            .I(N__2404));
    Span12Mux_v I__400 (
            .O(N__2407),
            .I(N__2401));
    Span4Mux_h I__399 (
            .O(N__2404),
            .I(N__2398));
    Odrv12 I__398 (
            .O(N__2401),
            .I(DIVIDE_8_));
    Odrv4 I__397 (
            .O(N__2398),
            .I(DIVIDE_8_));
    InMux I__396 (
            .O(N__2393),
            .I(N__2390));
    LocalMux I__395 (
            .O(N__2390),
            .I(t0on_15_N_35_7));
    CascadeMux I__394 (
            .O(N__2387),
            .I(N__2383));
    InMux I__393 (
            .O(N__2386),
            .I(N__2380));
    InMux I__392 (
            .O(N__2383),
            .I(N__2377));
    LocalMux I__391 (
            .O(N__2380),
            .I(t0on_7));
    LocalMux I__390 (
            .O(N__2377),
            .I(t0on_7));
    CascadeMux I__389 (
            .O(N__2372),
            .I(N__2368));
    InMux I__388 (
            .O(N__2371),
            .I(N__2365));
    InMux I__387 (
            .O(N__2368),
            .I(N__2362));
    LocalMux I__386 (
            .O(N__2365),
            .I(t0on_15));
    LocalMux I__385 (
            .O(N__2362),
            .I(t0on_15));
    InMux I__384 (
            .O(N__2357),
            .I(N__2354));
    LocalMux I__383 (
            .O(N__2354),
            .I(t0on_15_N_35_11));
    CascadeMux I__382 (
            .O(N__2351),
            .I(N__2348));
    InMux I__381 (
            .O(N__2348),
            .I(N__2345));
    LocalMux I__380 (
            .O(N__2345),
            .I(N__2341));
    InMux I__379 (
            .O(N__2344),
            .I(N__2338));
    Odrv4 I__378 (
            .O(N__2341),
            .I(t0on_11));
    LocalMux I__377 (
            .O(N__2338),
            .I(t0on_11));
    InMux I__376 (
            .O(N__2333),
            .I(n392));
    InMux I__375 (
            .O(N__2330),
            .I(n393));
    InMux I__374 (
            .O(N__2327),
            .I(n394));
    InMux I__373 (
            .O(N__2324),
            .I(bfn_2_10_0_));
    InMux I__372 (
            .O(N__2321),
            .I(n396));
    InMux I__371 (
            .O(N__2318),
            .I(n397));
    InMux I__370 (
            .O(N__2315),
            .I(n398));
    InMux I__369 (
            .O(N__2312),
            .I(n399));
    InMux I__368 (
            .O(N__2309),
            .I(n400));
    InMux I__367 (
            .O(N__2306),
            .I(n401));
    InMux I__366 (
            .O(N__2303),
            .I(n414));
    CascadeMux I__365 (
            .O(N__2300),
            .I(N__2297));
    InMux I__364 (
            .O(N__2297),
            .I(N__2293));
    InMux I__363 (
            .O(N__2296),
            .I(N__2290));
    LocalMux I__362 (
            .O(N__2293),
            .I(t0on_13));
    LocalMux I__361 (
            .O(N__2290),
            .I(t0on_13));
    InMux I__360 (
            .O(N__2285),
            .I(N__2282));
    LocalMux I__359 (
            .O(N__2282),
            .I(t0on_15_N_35_13));
    InMux I__358 (
            .O(N__2279),
            .I(n415));
    InMux I__357 (
            .O(N__2276),
            .I(n416));
    InMux I__356 (
            .O(N__2273),
            .I(n417));
    InMux I__355 (
            .O(N__2270),
            .I(bfn_2_9_0_));
    InMux I__354 (
            .O(N__2267),
            .I(n388));
    InMux I__353 (
            .O(N__2264),
            .I(n389));
    InMux I__352 (
            .O(N__2261),
            .I(n390));
    InMux I__351 (
            .O(N__2258),
            .I(n391));
    CascadeMux I__350 (
            .O(N__2255),
            .I(N__2251));
    InMux I__349 (
            .O(N__2254),
            .I(N__2248));
    InMux I__348 (
            .O(N__2251),
            .I(N__2245));
    LocalMux I__347 (
            .O(N__2248),
            .I(t0on_4));
    LocalMux I__346 (
            .O(N__2245),
            .I(t0on_4));
    InMux I__345 (
            .O(N__2240),
            .I(N__2237));
    LocalMux I__344 (
            .O(N__2237),
            .I(t0on_15_N_35_4));
    InMux I__343 (
            .O(N__2234),
            .I(n406));
    CascadeMux I__342 (
            .O(N__2231),
            .I(N__2227));
    CascadeMux I__341 (
            .O(N__2230),
            .I(N__2224));
    InMux I__340 (
            .O(N__2227),
            .I(N__2221));
    InMux I__339 (
            .O(N__2224),
            .I(N__2218));
    LocalMux I__338 (
            .O(N__2221),
            .I(t0on_5));
    LocalMux I__337 (
            .O(N__2218),
            .I(t0on_5));
    InMux I__336 (
            .O(N__2213),
            .I(N__2210));
    LocalMux I__335 (
            .O(N__2210),
            .I(t0on_15_N_35_5));
    InMux I__334 (
            .O(N__2207),
            .I(n407));
    InMux I__333 (
            .O(N__2204),
            .I(N__2200));
    InMux I__332 (
            .O(N__2203),
            .I(N__2197));
    LocalMux I__331 (
            .O(N__2200),
            .I(t0on_6));
    LocalMux I__330 (
            .O(N__2197),
            .I(t0on_6));
    InMux I__329 (
            .O(N__2192),
            .I(N__2189));
    LocalMux I__328 (
            .O(N__2189),
            .I(t0on_15_N_35_6));
    InMux I__327 (
            .O(N__2186),
            .I(n408));
    InMux I__326 (
            .O(N__2183),
            .I(n409));
    InMux I__325 (
            .O(N__2180),
            .I(N__2176));
    InMux I__324 (
            .O(N__2179),
            .I(N__2173));
    LocalMux I__323 (
            .O(N__2176),
            .I(t0on_8));
    LocalMux I__322 (
            .O(N__2173),
            .I(t0on_8));
    InMux I__321 (
            .O(N__2168),
            .I(N__2165));
    LocalMux I__320 (
            .O(N__2165),
            .I(t0on_15_N_35_8));
    InMux I__319 (
            .O(N__2162),
            .I(bfn_2_8_0_));
    InMux I__318 (
            .O(N__2159),
            .I(n411));
    InMux I__317 (
            .O(N__2156),
            .I(n412));
    InMux I__316 (
            .O(N__2153),
            .I(n413));
    InMux I__315 (
            .O(N__2150),
            .I(N__2147));
    LocalMux I__314 (
            .O(N__2147),
            .I(n3));
    InMux I__313 (
            .O(N__2144),
            .I(N__2140));
    CascadeMux I__312 (
            .O(N__2143),
            .I(N__2137));
    LocalMux I__311 (
            .O(N__2140),
            .I(N__2133));
    InMux I__310 (
            .O(N__2137),
            .I(N__2130));
    InMux I__309 (
            .O(N__2136),
            .I(N__2127));
    Span4Mux_v I__308 (
            .O(N__2133),
            .I(N__2122));
    LocalMux I__307 (
            .O(N__2130),
            .I(N__2122));
    LocalMux I__306 (
            .O(N__2127),
            .I(N__2119));
    Span4Mux_v I__305 (
            .O(N__2122),
            .I(N__2116));
    Span4Mux_v I__304 (
            .O(N__2119),
            .I(N__2113));
    Span4Mux_h I__303 (
            .O(N__2116),
            .I(N__2108));
    Span4Mux_h I__302 (
            .O(N__2113),
            .I(N__2108));
    Odrv4 I__301 (
            .O(N__2108),
            .I(DIVIDE_1_));
    InMux I__300 (
            .O(N__2105),
            .I(N__2102));
    LocalMux I__299 (
            .O(N__2102),
            .I(N__2099));
    Odrv4 I__298 (
            .O(N__2099),
            .I(n17));
    CascadeMux I__297 (
            .O(N__2096),
            .I(N__2093));
    InMux I__296 (
            .O(N__2093),
            .I(N__2090));
    LocalMux I__295 (
            .O(N__2090),
            .I(N__2086));
    InMux I__294 (
            .O(N__2089),
            .I(N__2083));
    Span4Mux_v I__293 (
            .O(N__2086),
            .I(N__2079));
    LocalMux I__292 (
            .O(N__2083),
            .I(N__2076));
    InMux I__291 (
            .O(N__2082),
            .I(N__2073));
    Span4Mux_h I__290 (
            .O(N__2079),
            .I(N__2070));
    Sp12to4 I__289 (
            .O(N__2076),
            .I(N__2065));
    LocalMux I__288 (
            .O(N__2073),
            .I(N__2065));
    Odrv4 I__287 (
            .O(N__2070),
            .I(DIVIDE_7_));
    Odrv12 I__286 (
            .O(N__2065),
            .I(DIVIDE_7_));
    CascadeMux I__285 (
            .O(N__2060),
            .I(N__2057));
    InMux I__284 (
            .O(N__2057),
            .I(N__2053));
    InMux I__283 (
            .O(N__2056),
            .I(N__2050));
    LocalMux I__282 (
            .O(N__2053),
            .I(N__2046));
    LocalMux I__281 (
            .O(N__2050),
            .I(N__2043));
    InMux I__280 (
            .O(N__2049),
            .I(N__2040));
    Sp12to4 I__279 (
            .O(N__2046),
            .I(N__2033));
    Sp12to4 I__278 (
            .O(N__2043),
            .I(N__2033));
    LocalMux I__277 (
            .O(N__2040),
            .I(N__2033));
    Span12Mux_v I__276 (
            .O(N__2033),
            .I(N__2030));
    Odrv12 I__275 (
            .O(N__2030),
            .I(DIVIDE_2_));
    InMux I__274 (
            .O(N__2027),
            .I(N__2023));
    InMux I__273 (
            .O(N__2026),
            .I(N__2020));
    LocalMux I__272 (
            .O(N__2023),
            .I(t0on_0));
    LocalMux I__271 (
            .O(N__2020),
            .I(t0on_0));
    InMux I__270 (
            .O(N__2015),
            .I(N__2012));
    LocalMux I__269 (
            .O(N__2012),
            .I(t0on_15_N_35_0));
    InMux I__268 (
            .O(N__2009),
            .I(bfn_2_7_0_));
    InMux I__267 (
            .O(N__2006),
            .I(N__2002));
    InMux I__266 (
            .O(N__2005),
            .I(N__1999));
    LocalMux I__265 (
            .O(N__2002),
            .I(t0on_1));
    LocalMux I__264 (
            .O(N__1999),
            .I(t0on_1));
    InMux I__263 (
            .O(N__1994),
            .I(N__1991));
    LocalMux I__262 (
            .O(N__1991),
            .I(t0on_15_N_35_1));
    InMux I__261 (
            .O(N__1988),
            .I(n403));
    InMux I__260 (
            .O(N__1985),
            .I(n404));
    InMux I__259 (
            .O(N__1982),
            .I(N__1978));
    InMux I__258 (
            .O(N__1981),
            .I(N__1975));
    LocalMux I__257 (
            .O(N__1978),
            .I(t0on_3));
    LocalMux I__256 (
            .O(N__1975),
            .I(t0on_3));
    InMux I__255 (
            .O(N__1970),
            .I(N__1967));
    LocalMux I__254 (
            .O(N__1967),
            .I(t0on_15_N_35_3));
    InMux I__253 (
            .O(N__1964),
            .I(n405));
    CascadeMux I__252 (
            .O(N__1961),
            .I(N__1958));
    InMux I__251 (
            .O(N__1958),
            .I(N__1955));
    LocalMux I__250 (
            .O(N__1955),
            .I(N__1952));
    Odrv4 I__249 (
            .O(N__1952),
            .I(n5));
    InMux I__248 (
            .O(N__1949),
            .I(n429));
    CascadeMux I__247 (
            .O(N__1946),
            .I(N__1943));
    InMux I__246 (
            .O(N__1943),
            .I(N__1940));
    LocalMux I__245 (
            .O(N__1940),
            .I(N__1937));
    Odrv4 I__244 (
            .O(N__1937),
            .I(n4));
    InMux I__243 (
            .O(N__1934),
            .I(n430));
    CascadeMux I__242 (
            .O(N__1931),
            .I(N__1928));
    InMux I__241 (
            .O(N__1928),
            .I(N__1923));
    InMux I__240 (
            .O(N__1927),
            .I(N__1920));
    InMux I__239 (
            .O(N__1926),
            .I(N__1917));
    LocalMux I__238 (
            .O(N__1923),
            .I(N__1910));
    LocalMux I__237 (
            .O(N__1920),
            .I(N__1910));
    LocalMux I__236 (
            .O(N__1917),
            .I(N__1910));
    Span4Mux_v I__235 (
            .O(N__1910),
            .I(N__1907));
    Span4Mux_v I__234 (
            .O(N__1907),
            .I(N__1904));
    Span4Mux_v I__233 (
            .O(N__1904),
            .I(N__1901));
    Sp12to4 I__232 (
            .O(N__1901),
            .I(N__1898));
    Odrv12 I__231 (
            .O(N__1898),
            .I(DIVIDE_14_));
    InMux I__230 (
            .O(N__1895),
            .I(n431));
    InMux I__229 (
            .O(N__1892),
            .I(n432));
    CascadeMux I__228 (
            .O(N__1889),
            .I(N__1886));
    InMux I__227 (
            .O(N__1886),
            .I(N__1883));
    LocalMux I__226 (
            .O(N__1883),
            .I(n7));
    IoInMux I__225 (
            .O(N__1880),
            .I(N__1877));
    LocalMux I__224 (
            .O(N__1877),
            .I(N__1874));
    Span12Mux_s4_h I__223 (
            .O(N__1874),
            .I(N__1871));
    Odrv12 I__222 (
            .O(N__1871),
            .I(OCLK));
    InMux I__221 (
            .O(N__1868),
            .I(N__1865));
    LocalMux I__220 (
            .O(N__1865),
            .I(N__1862));
    Odrv4 I__219 (
            .O(N__1862),
            .I(n10));
    InMux I__218 (
            .O(N__1859),
            .I(N__1855));
    InMux I__217 (
            .O(N__1858),
            .I(N__1852));
    LocalMux I__216 (
            .O(N__1855),
            .I(N__1846));
    LocalMux I__215 (
            .O(N__1852),
            .I(N__1846));
    InMux I__214 (
            .O(N__1851),
            .I(N__1843));
    Span4Mux_v I__213 (
            .O(N__1846),
            .I(N__1838));
    LocalMux I__212 (
            .O(N__1843),
            .I(N__1838));
    Span4Mux_v I__211 (
            .O(N__1838),
            .I(N__1835));
    Span4Mux_h I__210 (
            .O(N__1835),
            .I(N__1832));
    Odrv4 I__209 (
            .O(N__1832),
            .I(DIVIDE_6_));
    InMux I__208 (
            .O(N__1829),
            .I(N__1826));
    LocalMux I__207 (
            .O(N__1826),
            .I(N__1823));
    Odrv4 I__206 (
            .O(N__1823),
            .I(n12));
    InMux I__205 (
            .O(N__1820),
            .I(N__1817));
    LocalMux I__204 (
            .O(N__1817),
            .I(n14));
    InMux I__203 (
            .O(N__1814),
            .I(n420));
    InMux I__202 (
            .O(N__1811),
            .I(N__1808));
    LocalMux I__201 (
            .O(N__1808),
            .I(n13));
    CascadeMux I__200 (
            .O(N__1805),
            .I(N__1802));
    InMux I__199 (
            .O(N__1802),
            .I(N__1799));
    LocalMux I__198 (
            .O(N__1799),
            .I(N__1794));
    InMux I__197 (
            .O(N__1798),
            .I(N__1791));
    InMux I__196 (
            .O(N__1797),
            .I(N__1788));
    Span4Mux_v I__195 (
            .O(N__1794),
            .I(N__1781));
    LocalMux I__194 (
            .O(N__1791),
            .I(N__1781));
    LocalMux I__193 (
            .O(N__1788),
            .I(N__1781));
    Span4Mux_v I__192 (
            .O(N__1781),
            .I(N__1778));
    Span4Mux_h I__191 (
            .O(N__1778),
            .I(N__1775));
    Span4Mux_v I__190 (
            .O(N__1775),
            .I(N__1772));
    Odrv4 I__189 (
            .O(N__1772),
            .I(DIVIDE_4_));
    InMux I__188 (
            .O(N__1769),
            .I(n421));
    CascadeMux I__187 (
            .O(N__1766),
            .I(N__1763));
    InMux I__186 (
            .O(N__1763),
            .I(N__1759));
    InMux I__185 (
            .O(N__1762),
            .I(N__1756));
    LocalMux I__184 (
            .O(N__1759),
            .I(N__1751));
    LocalMux I__183 (
            .O(N__1756),
            .I(N__1751));
    Span4Mux_v I__182 (
            .O(N__1751),
            .I(N__1747));
    InMux I__181 (
            .O(N__1750),
            .I(N__1744));
    Sp12to4 I__180 (
            .O(N__1747),
            .I(N__1739));
    LocalMux I__179 (
            .O(N__1744),
            .I(N__1739));
    Odrv12 I__178 (
            .O(N__1739),
            .I(DIVIDE_5_));
    InMux I__177 (
            .O(N__1736),
            .I(n422));
    CascadeMux I__176 (
            .O(N__1733),
            .I(N__1730));
    InMux I__175 (
            .O(N__1730),
            .I(N__1727));
    LocalMux I__174 (
            .O(N__1727),
            .I(N__1724));
    Odrv4 I__173 (
            .O(N__1724),
            .I(n11));
    InMux I__172 (
            .O(N__1721),
            .I(n423));
    InMux I__171 (
            .O(N__1718),
            .I(n424));
    CascadeMux I__170 (
            .O(N__1715),
            .I(N__1712));
    InMux I__169 (
            .O(N__1712),
            .I(N__1709));
    LocalMux I__168 (
            .O(N__1709),
            .I(N__1706));
    Odrv4 I__167 (
            .O(N__1706),
            .I(n9));
    InMux I__166 (
            .O(N__1703),
            .I(bfn_1_10_0_));
    InMux I__165 (
            .O(N__1700),
            .I(N__1695));
    InMux I__164 (
            .O(N__1699),
            .I(N__1692));
    InMux I__163 (
            .O(N__1698),
            .I(N__1689));
    LocalMux I__162 (
            .O(N__1695),
            .I(N__1686));
    LocalMux I__161 (
            .O(N__1692),
            .I(N__1681));
    LocalMux I__160 (
            .O(N__1689),
            .I(N__1681));
    Sp12to4 I__159 (
            .O(N__1686),
            .I(N__1678));
    Span4Mux_v I__158 (
            .O(N__1681),
            .I(N__1675));
    Span12Mux_s5_h I__157 (
            .O(N__1678),
            .I(N__1670));
    Sp12to4 I__156 (
            .O(N__1675),
            .I(N__1670));
    Span12Mux_v I__155 (
            .O(N__1670),
            .I(N__1667));
    Odrv12 I__154 (
            .O(N__1667),
            .I(DIVIDE_9_));
    InMux I__153 (
            .O(N__1664),
            .I(n426));
    InMux I__152 (
            .O(N__1661),
            .I(n427));
    InMux I__151 (
            .O(N__1658),
            .I(n428));
    CascadeMux I__150 (
            .O(N__1655),
            .I(N__1652));
    InMux I__149 (
            .O(N__1652),
            .I(N__1649));
    LocalMux I__148 (
            .O(N__1649),
            .I(N__1646));
    Sp12to4 I__147 (
            .O(N__1646),
            .I(N__1643));
    Span12Mux_v I__146 (
            .O(N__1643),
            .I(N__1640));
    Odrv12 I__145 (
            .O(N__1640),
            .I(DIVIDE_0_));
    InMux I__144 (
            .O(N__1637),
            .I(bfn_1_9_0_));
    InMux I__143 (
            .O(N__1634),
            .I(N__1631));
    LocalMux I__142 (
            .O(N__1631),
            .I(n16));
    InMux I__141 (
            .O(N__1628),
            .I(n418));
    InMux I__140 (
            .O(N__1625),
            .I(N__1622));
    LocalMux I__139 (
            .O(N__1622),
            .I(n15));
    InMux I__138 (
            .O(N__1619),
            .I(n419));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(n425),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(n395),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(n410),
            .carryinitout(bfn_2_8_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i200_4_lut_LC_1_6_0.C_ON=1'b0;
    defparam i200_4_lut_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam i200_4_lut_LC_1_6_0.LUT_INIT=16'b1111111111111011;
    LogicCell40 i200_4_lut_LC_1_6_0 (
            .in0(N__2203),
            .in1(N__2005),
            .in2(N__2255),
            .in3(N__2026),
            .lcout(n447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i4_LC_1_6_3.C_ON=1'b0;
    defparam t0on_i4_LC_1_6_3.SEQ_MODE=4'b1000;
    defparam t0on_i4_LC_1_6_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0on_i4_LC_1_6_3 (
            .in0(N__1750),
            .in1(N__3344),
            .in2(_gnd_net_),
            .in3(N__2240),
            .lcout(t0on_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3678),
            .ce(N__3406),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i7_1_lut_LC_1_6_5.C_ON=1'b0;
    defparam sub_34_inv_0_i7_1_lut_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i7_1_lut_LC_1_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i7_1_lut_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2082),
            .lcout(n11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i0_LC_1_7_0.C_ON=1'b0;
    defparam t0on_i0_LC_1_7_0.SEQ_MODE=4'b1000;
    defparam t0on_i0_LC_1_7_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0on_i0_LC_1_7_0 (
            .in0(N__2144),
            .in1(N__3337),
            .in2(_gnd_net_),
            .in3(N__2015),
            .lcout(t0on_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3680),
            .ce(N__3412),
            .sr(_gnd_net_));
    defparam t0on_i8_LC_1_7_1.C_ON=1'b0;
    defparam t0on_i8_LC_1_7_1.SEQ_MODE=4'b1000;
    defparam t0on_i8_LC_1_7_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i8_LC_1_7_1 (
            .in0(N__3341),
            .in1(N__1698),
            .in2(_gnd_net_),
            .in3(N__2168),
            .lcout(t0on_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3680),
            .ce(N__3412),
            .sr(_gnd_net_));
    defparam t0on_i13_LC_1_7_5.C_ON=1'b0;
    defparam t0on_i13_LC_1_7_5.SEQ_MODE=4'b1000;
    defparam t0on_i13_LC_1_7_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i13_LC_1_7_5 (
            .in0(N__3338),
            .in1(N__1926),
            .in2(_gnd_net_),
            .in3(N__2285),
            .lcout(t0on_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3680),
            .ce(N__3412),
            .sr(_gnd_net_));
    defparam t0on_i5_LC_1_7_6.C_ON=1'b0;
    defparam t0on_i5_LC_1_7_6.SEQ_MODE=4'b1000;
    defparam t0on_i5_LC_1_7_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0on_i5_LC_1_7_6 (
            .in0(N__1859),
            .in1(N__3340),
            .in2(_gnd_net_),
            .in3(N__2213),
            .lcout(t0on_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3680),
            .ce(N__3412),
            .sr(_gnd_net_));
    defparam t0on_i3_LC_1_7_7.C_ON=1'b0;
    defparam t0on_i3_LC_1_7_7.SEQ_MODE=4'b1000;
    defparam t0on_i3_LC_1_7_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i3_LC_1_7_7 (
            .in0(N__3339),
            .in1(N__1797),
            .in2(_gnd_net_),
            .in3(N__1970),
            .lcout(t0on_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3680),
            .ce(N__3412),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i2_1_lut_LC_1_8_0.C_ON=1'b0;
    defparam sub_34_inv_0_i2_1_lut_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i2_1_lut_LC_1_8_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i2_1_lut_LC_1_8_0 (
            .in0(N__2056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i5_1_lut_LC_1_8_1.C_ON=1'b0;
    defparam sub_34_inv_0_i5_1_lut_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i5_1_lut_LC_1_8_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i5_1_lut_LC_1_8_1 (
            .in0(N__1762),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i13_1_lut_LC_1_8_2.C_ON=1'b0;
    defparam sub_34_inv_0_i13_1_lut_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i13_1_lut_LC_1_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i13_1_lut_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2491),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i14_1_lut_LC_1_8_3.C_ON=1'b0;
    defparam sub_34_inv_0_i14_1_lut_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i14_1_lut_LC_1_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i14_1_lut_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1927),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i4_1_lut_LC_1_8_4.C_ON=1'b0;
    defparam sub_34_inv_0_i4_1_lut_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i4_1_lut_LC_1_8_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i4_1_lut_LC_1_8_4 (
            .in0(N__1798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_1_LC_1_8_5.C_ON=1'b0;
    defparam i10_4_lut_adj_1_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_1_LC_1_8_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_1_LC_1_8_5 (
            .in0(N__2296),
            .in1(N__1981),
            .in2(N__2230),
            .in3(N__2179),
            .lcout(n26_adj_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i9_1_lut_LC_1_8_6.C_ON=1'b0;
    defparam sub_34_inv_0_i9_1_lut_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i9_1_lut_LC_1_8_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i9_1_lut_LC_1_8_6 (
            .in0(N__1699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i3_1_lut_LC_1_8_7.C_ON=1'b0;
    defparam sub_34_inv_0_i3_1_lut_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i3_1_lut_LC_1_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i3_1_lut_LC_1_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2544),
            .lcout(n15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_2_lut_LC_1_9_0.C_ON=1'b1;
    defparam sub_34_add_2_2_lut_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_2_lut_LC_1_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_2_lut_LC_1_9_0 (
            .in0(_gnd_net_),
            .in1(N__2105),
            .in2(N__1655),
            .in3(N__1637),
            .lcout(t0off_15_N_67_0),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(n418),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_3_lut_LC_1_9_1.C_ON=1'b1;
    defparam sub_34_add_2_3_lut_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_3_lut_LC_1_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_3_lut_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(N__1634),
            .in2(N__2143),
            .in3(N__1628),
            .lcout(t0off_15_N_67_1),
            .ltout(),
            .carryin(n418),
            .carryout(n419),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_4_lut_LC_1_9_2.C_ON=1'b1;
    defparam sub_34_add_2_4_lut_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_4_lut_LC_1_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_4_lut_LC_1_9_2 (
            .in0(_gnd_net_),
            .in1(N__1625),
            .in2(N__2060),
            .in3(N__1619),
            .lcout(t0off_15_N_67_2),
            .ltout(),
            .carryin(n419),
            .carryout(n420),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_5_lut_LC_1_9_3.C_ON=1'b1;
    defparam sub_34_add_2_5_lut_LC_1_9_3.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_5_lut_LC_1_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_5_lut_LC_1_9_3 (
            .in0(_gnd_net_),
            .in1(N__1820),
            .in2(N__2549),
            .in3(N__1814),
            .lcout(t0off_15_N_67_3),
            .ltout(),
            .carryin(n420),
            .carryout(n421),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_6_lut_LC_1_9_4.C_ON=1'b1;
    defparam sub_34_add_2_6_lut_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_6_lut_LC_1_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_6_lut_LC_1_9_4 (
            .in0(_gnd_net_),
            .in1(N__1811),
            .in2(N__1805),
            .in3(N__1769),
            .lcout(t0off_15_N_67_4),
            .ltout(),
            .carryin(n421),
            .carryout(n422),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_7_lut_LC_1_9_5.C_ON=1'b1;
    defparam sub_34_add_2_7_lut_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_7_lut_LC_1_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_7_lut_LC_1_9_5 (
            .in0(_gnd_net_),
            .in1(N__1829),
            .in2(N__1766),
            .in3(N__1736),
            .lcout(t0off_15_N_67_5),
            .ltout(),
            .carryin(n422),
            .carryout(n423),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_8_lut_LC_1_9_6.C_ON=1'b1;
    defparam sub_34_add_2_8_lut_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_8_lut_LC_1_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_8_lut_LC_1_9_6 (
            .in0(_gnd_net_),
            .in1(N__1858),
            .in2(N__1733),
            .in3(N__1721),
            .lcout(t0off_15_N_67_6),
            .ltout(),
            .carryin(n423),
            .carryout(n424),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_9_lut_LC_1_9_7.C_ON=1'b1;
    defparam sub_34_add_2_9_lut_LC_1_9_7.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_9_lut_LC_1_9_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_9_lut_LC_1_9_7 (
            .in0(_gnd_net_),
            .in1(N__1868),
            .in2(N__2096),
            .in3(N__1718),
            .lcout(t0off_15_N_67_7),
            .ltout(),
            .carryin(n424),
            .carryout(n425),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_10_lut_LC_1_10_0.C_ON=1'b1;
    defparam sub_34_add_2_10_lut_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_10_lut_LC_1_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_10_lut_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(N__2434),
            .in2(N__1715),
            .in3(N__1703),
            .lcout(t0off_15_N_67_8),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(n426),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_11_lut_LC_1_10_1.C_ON=1'b1;
    defparam sub_34_add_2_11_lut_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_11_lut_LC_1_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_11_lut_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(N__1700),
            .in2(N__2894),
            .in3(N__1664),
            .lcout(t0off_15_N_67_9),
            .ltout(),
            .carryin(n426),
            .carryout(n427),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_12_lut_LC_1_10_2.C_ON=1'b1;
    defparam sub_34_add_2_12_lut_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_12_lut_LC_1_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_12_lut_LC_1_10_2 (
            .in0(_gnd_net_),
            .in1(N__2908),
            .in2(N__1889),
            .in3(N__1661),
            .lcout(t0off_15_N_67_10),
            .ltout(),
            .carryin(n427),
            .carryout(n428),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_13_lut_LC_1_10_3.C_ON=1'b1;
    defparam sub_34_add_2_13_lut_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_13_lut_LC_1_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_13_lut_LC_1_10_3 (
            .in0(_gnd_net_),
            .in1(N__2930),
            .in2(N__2609),
            .in3(N__1658),
            .lcout(t0off_15_N_67_11),
            .ltout(),
            .carryin(n428),
            .carryout(n429),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_14_lut_LC_1_10_4.C_ON=1'b1;
    defparam sub_34_add_2_14_lut_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_14_lut_LC_1_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_14_lut_LC_1_10_4 (
            .in0(_gnd_net_),
            .in1(N__2944),
            .in2(N__1961),
            .in3(N__1949),
            .lcout(t0off_15_N_67_12),
            .ltout(),
            .carryin(n429),
            .carryout(n430),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_15_lut_LC_1_10_5.C_ON=1'b1;
    defparam sub_34_add_2_15_lut_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_15_lut_LC_1_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_15_lut_LC_1_10_5 (
            .in0(_gnd_net_),
            .in1(N__2495),
            .in2(N__1946),
            .in3(N__1934),
            .lcout(t0off_15_N_67_13),
            .ltout(),
            .carryin(n430),
            .carryout(n431),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_add_2_16_lut_LC_1_10_6.C_ON=1'b1;
    defparam sub_34_add_2_16_lut_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam sub_34_add_2_16_lut_LC_1_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sub_34_add_2_16_lut_LC_1_10_6 (
            .in0(_gnd_net_),
            .in1(N__2150),
            .in2(N__1931),
            .in3(N__1895),
            .lcout(t0off_15_N_67_14),
            .ltout(),
            .carryin(n431),
            .carryout(n432),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0off_i15_LC_1_10_7.C_ON=1'b0;
    defparam t0off_i15_LC_1_10_7.SEQ_MODE=4'b1000;
    defparam t0off_i15_LC_1_10_7.LUT_INIT=16'b1011100001110100;
    LogicCell40 t0off_i15_LC_1_10_7 (
            .in0(N__3007),
            .in1(N__3402),
            .in2(N__2618),
            .in3(N__1892),
            .lcout(t0off_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3648),
            .ce(N__3545),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i11_1_lut_LC_1_11_0.C_ON=1'b0;
    defparam sub_34_inv_0_i11_1_lut_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i11_1_lut_LC_1_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i11_1_lut_LC_1_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2607),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t_clk_24_LC_1_11_1.C_ON=1'b0;
    defparam t_clk_24_LC_1_11_1.SEQ_MODE=4'b1000;
    defparam t_clk_24_LC_1_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 t_clk_24_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3811),
            .lcout(OCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3614),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i8_1_lut_LC_1_11_2.C_ON=1'b0;
    defparam sub_34_inv_0_i8_1_lut_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i8_1_lut_LC_1_11_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i8_1_lut_LC_1_11_2 (
            .in0(N__2433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i6_1_lut_LC_1_11_4.C_ON=1'b0;
    defparam sub_34_inv_0_i6_1_lut_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i6_1_lut_LC_1_11_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 sub_34_inv_0_i6_1_lut_LC_1_11_4 (
            .in0(N__1851),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i15_1_lut_LC_1_11_5.C_ON=1'b0;
    defparam sub_34_inv_0_i15_1_lut_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i15_1_lut_LC_1_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i15_1_lut_LC_1_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2994),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i1_1_lut_LC_1_11_7.C_ON=1'b0;
    defparam sub_34_inv_0_i1_1_lut_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i1_1_lut_LC_1_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i1_1_lut_LC_1_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2136),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_5_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_5_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_5_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i6_LC_2_6_5.C_ON=1'b0;
    defparam t0on_i6_LC_2_6_5.SEQ_MODE=4'b1000;
    defparam t0on_i6_LC_2_6_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i6_LC_2_6_5 (
            .in0(N__3343),
            .in1(N__2089),
            .in2(_gnd_net_),
            .in3(N__2192),
            .lcout(t0on_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3679),
            .ce(N__3407),
            .sr(_gnd_net_));
    defparam t0on_i1_LC_2_6_6.C_ON=1'b0;
    defparam t0on_i1_LC_2_6_6.SEQ_MODE=4'b1000;
    defparam t0on_i1_LC_2_6_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 t0on_i1_LC_2_6_6 (
            .in0(N__2049),
            .in1(N__1994),
            .in2(_gnd_net_),
            .in3(N__3342),
            .lcout(t0on_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3679),
            .ce(N__3407),
            .sr(_gnd_net_));
    defparam add_32_2_lut_LC_2_7_0.C_ON=1'b1;
    defparam add_32_2_lut_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam add_32_2_lut_LC_2_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_2_lut_LC_2_7_0 (
            .in0(_gnd_net_),
            .in1(N__2027),
            .in2(_gnd_net_),
            .in3(N__2009),
            .lcout(t0on_15_N_35_0),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(n403),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_3_lut_LC_2_7_1.C_ON=1'b1;
    defparam add_32_3_lut_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam add_32_3_lut_LC_2_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_3_lut_LC_2_7_1 (
            .in0(_gnd_net_),
            .in1(N__2006),
            .in2(N__2768),
            .in3(N__1988),
            .lcout(t0on_15_N_35_1),
            .ltout(),
            .carryin(n403),
            .carryout(n404),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_4_lut_LC_2_7_2.C_ON=1'b1;
    defparam add_32_4_lut_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam add_32_4_lut_LC_2_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_4_lut_LC_2_7_2 (
            .in0(_gnd_net_),
            .in1(N__2507),
            .in2(N__2771),
            .in3(N__1985),
            .lcout(t0on_15_N_35_2),
            .ltout(),
            .carryin(n404),
            .carryout(n405),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_5_lut_LC_2_7_3.C_ON=1'b1;
    defparam add_32_5_lut_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam add_32_5_lut_LC_2_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_5_lut_LC_2_7_3 (
            .in0(_gnd_net_),
            .in1(N__1982),
            .in2(N__2769),
            .in3(N__1964),
            .lcout(t0on_15_N_35_3),
            .ltout(),
            .carryin(n405),
            .carryout(n406),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_6_lut_LC_2_7_4.C_ON=1'b1;
    defparam add_32_6_lut_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam add_32_6_lut_LC_2_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_6_lut_LC_2_7_4 (
            .in0(_gnd_net_),
            .in1(N__2254),
            .in2(N__2772),
            .in3(N__2234),
            .lcout(t0on_15_N_35_4),
            .ltout(),
            .carryin(n406),
            .carryout(n407),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_7_lut_LC_2_7_5.C_ON=1'b1;
    defparam add_32_7_lut_LC_2_7_5.SEQ_MODE=4'b0000;
    defparam add_32_7_lut_LC_2_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_7_lut_LC_2_7_5 (
            .in0(_gnd_net_),
            .in1(N__2709),
            .in2(N__2231),
            .in3(N__2207),
            .lcout(t0on_15_N_35_5),
            .ltout(),
            .carryin(n407),
            .carryout(n408),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_8_lut_LC_2_7_6.C_ON=1'b1;
    defparam add_32_8_lut_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam add_32_8_lut_LC_2_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_8_lut_LC_2_7_6 (
            .in0(_gnd_net_),
            .in1(N__2204),
            .in2(N__2773),
            .in3(N__2186),
            .lcout(t0on_15_N_35_6),
            .ltout(),
            .carryin(n408),
            .carryout(n409),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_9_lut_LC_2_7_7.C_ON=1'b1;
    defparam add_32_9_lut_LC_2_7_7.SEQ_MODE=4'b0000;
    defparam add_32_9_lut_LC_2_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_9_lut_LC_2_7_7 (
            .in0(_gnd_net_),
            .in1(N__2386),
            .in2(N__2770),
            .in3(N__2183),
            .lcout(t0on_15_N_35_7),
            .ltout(),
            .carryin(n409),
            .carryout(n410),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_10_lut_LC_2_8_0.C_ON=1'b1;
    defparam add_32_10_lut_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam add_32_10_lut_LC_2_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_10_lut_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(N__2180),
            .in2(N__2774),
            .in3(N__2162),
            .lcout(t0on_15_N_35_8),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(n411),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_11_lut_LC_2_8_1.C_ON=1'b1;
    defparam add_32_11_lut_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam add_32_11_lut_LC_2_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_11_lut_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(N__2716),
            .in2(N__3023),
            .in3(N__2159),
            .lcout(t0on_15_N_35_9),
            .ltout(),
            .carryin(n411),
            .carryout(n412),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_12_lut_LC_2_8_2.C_ON=1'b1;
    defparam add_32_12_lut_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam add_32_12_lut_LC_2_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_12_lut_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(N__2561),
            .in2(N__2775),
            .in3(N__2156),
            .lcout(t0on_15_N_35_10),
            .ltout(),
            .carryin(n412),
            .carryout(n413),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_13_lut_LC_2_8_3.C_ON=1'b1;
    defparam add_32_13_lut_LC_2_8_3.SEQ_MODE=4'b0000;
    defparam add_32_13_lut_LC_2_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_13_lut_LC_2_8_3 (
            .in0(_gnd_net_),
            .in1(N__2720),
            .in2(N__2351),
            .in3(N__2153),
            .lcout(t0on_15_N_35_11),
            .ltout(),
            .carryin(n413),
            .carryout(n414),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_14_lut_LC_2_8_4.C_ON=1'b1;
    defparam add_32_14_lut_LC_2_8_4.SEQ_MODE=4'b0000;
    defparam add_32_14_lut_LC_2_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_14_lut_LC_2_8_4 (
            .in0(_gnd_net_),
            .in1(N__2447),
            .in2(N__2776),
            .in3(N__2303),
            .lcout(t0on_15_N_35_12),
            .ltout(),
            .carryin(n414),
            .carryout(n415),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_15_lut_LC_2_8_5.C_ON=1'b1;
    defparam add_32_15_lut_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam add_32_15_lut_LC_2_8_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_15_lut_LC_2_8_5 (
            .in0(_gnd_net_),
            .in1(N__2724),
            .in2(N__2300),
            .in3(N__2279),
            .lcout(t0on_15_N_35_13),
            .ltout(),
            .carryin(n415),
            .carryout(n416),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_32_16_lut_LC_2_8_6.C_ON=1'b1;
    defparam add_32_16_lut_LC_2_8_6.SEQ_MODE=4'b0000;
    defparam add_32_16_lut_LC_2_8_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_32_16_lut_LC_2_8_6 (
            .in0(_gnd_net_),
            .in1(N__2969),
            .in2(N__2777),
            .in3(N__2276),
            .lcout(t0on_15_N_35_14),
            .ltout(),
            .carryin(n416),
            .carryout(n417),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i15_LC_2_8_7.C_ON=1'b0;
    defparam t0on_i15_LC_2_8_7.SEQ_MODE=4'b1000;
    defparam t0on_i15_LC_2_8_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 t0on_i15_LC_2_8_7 (
            .in0(N__2371),
            .in1(N__2728),
            .in2(_gnd_net_),
            .in3(N__2273),
            .lcout(t0on_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3681),
            .ce(N__3413),
            .sr(N__3425));
    defparam add_33_2_lut_LC_2_9_0.C_ON=1'b1;
    defparam add_33_2_lut_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam add_33_2_lut_LC_2_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_2_lut_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(N__3931),
            .in2(_gnd_net_),
            .in3(N__2270),
            .lcout(t0off_15_N_51_0),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(n388),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_3_lut_LC_2_9_1.C_ON=1'b1;
    defparam add_33_3_lut_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam add_33_3_lut_LC_2_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_3_lut_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__3964),
            .in2(N__2778),
            .in3(N__2267),
            .lcout(t0off_15_N_51_1),
            .ltout(),
            .carryin(n388),
            .carryout(n389),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_4_lut_LC_2_9_2.C_ON=1'b1;
    defparam add_33_4_lut_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam add_33_4_lut_LC_2_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_4_lut_LC_2_9_2 (
            .in0(_gnd_net_),
            .in1(N__3220),
            .in2(N__2782),
            .in3(N__2264),
            .lcout(t0off_15_N_51_2),
            .ltout(),
            .carryin(n389),
            .carryout(n390),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_5_lut_LC_2_9_3.C_ON=1'b1;
    defparam add_33_5_lut_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam add_33_5_lut_LC_2_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_5_lut_LC_2_9_3 (
            .in0(_gnd_net_),
            .in1(N__4055),
            .in2(N__2779),
            .in3(N__2261),
            .lcout(t0off_15_N_51_3),
            .ltout(),
            .carryin(n390),
            .carryout(n391),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_6_lut_LC_2_9_4.C_ON=1'b1;
    defparam add_33_6_lut_LC_2_9_4.SEQ_MODE=4'b0000;
    defparam add_33_6_lut_LC_2_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_6_lut_LC_2_9_4 (
            .in0(_gnd_net_),
            .in1(N__3946),
            .in2(N__2783),
            .in3(N__2258),
            .lcout(t0off_15_N_51_4),
            .ltout(),
            .carryin(n391),
            .carryout(n392),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_7_lut_LC_2_9_5.C_ON=1'b1;
    defparam add_33_7_lut_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam add_33_7_lut_LC_2_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_7_lut_LC_2_9_5 (
            .in0(_gnd_net_),
            .in1(N__3890),
            .in2(N__2780),
            .in3(N__2333),
            .lcout(t0off_15_N_51_5),
            .ltout(),
            .carryin(n392),
            .carryout(n393),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_8_lut_LC_2_9_6.C_ON=1'b1;
    defparam add_33_8_lut_LC_2_9_6.SEQ_MODE=4'b0000;
    defparam add_33_8_lut_LC_2_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_8_lut_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(N__3851),
            .in2(N__2784),
            .in3(N__2330),
            .lcout(t0off_15_N_51_6),
            .ltout(),
            .carryin(n393),
            .carryout(n394),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_9_lut_LC_2_9_7.C_ON=1'b1;
    defparam add_33_9_lut_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam add_33_9_lut_LC_2_9_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_9_lut_LC_2_9_7 (
            .in0(_gnd_net_),
            .in1(N__3202),
            .in2(N__2781),
            .in3(N__2327),
            .lcout(t0off_15_N_51_7),
            .ltout(),
            .carryin(n394),
            .carryout(n395),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_10_lut_LC_2_10_0.C_ON=1'b1;
    defparam add_33_10_lut_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam add_33_10_lut_LC_2_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_10_lut_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(N__4039),
            .in2(N__2805),
            .in3(N__2324),
            .lcout(t0off_15_N_51_8),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(n396),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_11_lut_LC_2_10_1.C_ON=1'b1;
    defparam add_33_11_lut_LC_2_10_1.SEQ_MODE=4'b0000;
    defparam add_33_11_lut_LC_2_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_11_lut_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(N__3986),
            .in2(N__2809),
            .in3(N__2321),
            .lcout(t0off_15_N_51_9),
            .ltout(),
            .carryin(n396),
            .carryout(n397),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_12_lut_LC_2_10_2.C_ON=1'b1;
    defparam add_33_12_lut_LC_2_10_2.SEQ_MODE=4'b0000;
    defparam add_33_12_lut_LC_2_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_12_lut_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(N__3187),
            .in2(N__2806),
            .in3(N__2318),
            .lcout(t0off_15_N_51_10),
            .ltout(),
            .carryin(n397),
            .carryout(n398),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_13_lut_LC_2_10_3.C_ON=1'b1;
    defparam add_33_13_lut_LC_2_10_3.SEQ_MODE=4'b0000;
    defparam add_33_13_lut_LC_2_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_13_lut_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(N__3707),
            .in2(N__2810),
            .in3(N__2315),
            .lcout(t0off_15_N_51_11),
            .ltout(),
            .carryin(n398),
            .carryout(n399),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_14_lut_LC_2_10_4.C_ON=1'b1;
    defparam add_33_14_lut_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam add_33_14_lut_LC_2_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_14_lut_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__3235),
            .in2(N__2807),
            .in3(N__2312),
            .lcout(t0off_15_N_51_12),
            .ltout(),
            .carryin(n399),
            .carryout(n400),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_15_lut_LC_2_10_5.C_ON=1'b1;
    defparam add_33_15_lut_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam add_33_15_lut_LC_2_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_15_lut_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(N__2794),
            .in2(N__4073),
            .in3(N__2309),
            .lcout(t0off_15_N_51_13),
            .ltout(),
            .carryin(n400),
            .carryout(n401),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_16_lut_LC_2_10_6.C_ON=1'b1;
    defparam add_33_16_lut_LC_2_10_6.SEQ_MODE=4'b0000;
    defparam add_33_16_lut_LC_2_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_33_16_lut_LC_2_10_6 (
            .in0(_gnd_net_),
            .in1(N__4018),
            .in2(N__2808),
            .in3(N__2306),
            .lcout(t0off_15_N_51_14),
            .ltout(),
            .carryin(n401),
            .carryout(n402),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_33_17_lut_LC_2_10_7.C_ON=1'b0;
    defparam add_33_17_lut_LC_2_10_7.SEQ_MODE=4'b0000;
    defparam add_33_17_lut_LC_2_10_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 add_33_17_lut_LC_2_10_7 (
            .in0(N__2804),
            .in1(N__4000),
            .in2(_gnd_net_),
            .in3(N__2621),
            .lcout(t0off_15_N_51_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_2_LC_3_7_0.C_ON=1'b0;
    defparam i11_4_lut_adj_2_LC_3_7_0.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_2_LC_3_7_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_2_LC_3_7_0 (
            .in0(N__2446),
            .in1(N__2506),
            .in2(N__2387),
            .in3(N__2560),
            .lcout(n27_adj_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i10_LC_3_7_1.C_ON=1'b0;
    defparam t0on_i10_LC_3_7_1.SEQ_MODE=4'b1000;
    defparam t0on_i10_LC_3_7_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0on_i10_LC_3_7_1 (
            .in0(N__2608),
            .in1(N__3333),
            .in2(_gnd_net_),
            .in3(N__2567),
            .lcout(t0on_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3691),
            .ce(N__3411),
            .sr(_gnd_net_));
    defparam t0on_i2_LC_3_7_2.C_ON=1'b0;
    defparam t0on_i2_LC_3_7_2.SEQ_MODE=4'b1000;
    defparam t0on_i2_LC_3_7_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i2_LC_3_7_2 (
            .in0(N__3335),
            .in1(N__2548),
            .in2(_gnd_net_),
            .in3(N__2513),
            .lcout(t0on_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3691),
            .ce(N__3411),
            .sr(_gnd_net_));
    defparam t0on_i12_LC_3_7_3.C_ON=1'b0;
    defparam t0on_i12_LC_3_7_3.SEQ_MODE=4'b1000;
    defparam t0on_i12_LC_3_7_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0on_i12_LC_3_7_3 (
            .in0(N__2490),
            .in1(N__3334),
            .in2(_gnd_net_),
            .in3(N__2453),
            .lcout(t0on_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3691),
            .ce(N__3411),
            .sr(_gnd_net_));
    defparam t0on_i7_LC_3_7_4.C_ON=1'b0;
    defparam t0on_i7_LC_3_7_4.SEQ_MODE=4'b1000;
    defparam t0on_i7_LC_3_7_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i7_LC_3_7_4 (
            .in0(N__3336),
            .in1(N__2435),
            .in2(_gnd_net_),
            .in3(N__2393),
            .lcout(t0on_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3691),
            .ce(N__3411),
            .sr(_gnd_net_));
    defparam i12_4_lut_LC_3_8_0.C_ON=1'b0;
    defparam i12_4_lut_LC_3_8_0.SEQ_MODE=4'b0000;
    defparam i12_4_lut_LC_3_8_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_LC_3_8_0 (
            .in0(N__2968),
            .in1(N__3019),
            .in2(N__2372),
            .in3(N__2344),
            .lcout(n28_adj_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0on_i11_LC_3_8_1.C_ON=1'b0;
    defparam t0on_i11_LC_3_8_1.SEQ_MODE=4'b1000;
    defparam t0on_i11_LC_3_8_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 t0on_i11_LC_3_8_1 (
            .in0(N__2357),
            .in1(_gnd_net_),
            .in2(N__3324),
            .in3(N__2957),
            .lcout(t0on_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3676),
            .ce(N__3398),
            .sr(_gnd_net_));
    defparam t0on_i9_LC_3_8_2.C_ON=1'b0;
    defparam t0on_i9_LC_3_8_2.SEQ_MODE=4'b1000;
    defparam t0on_i9_LC_3_8_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 t0on_i9_LC_3_8_2 (
            .in0(N__2918),
            .in1(N__3029),
            .in2(_gnd_net_),
            .in3(N__3298),
            .lcout(t0on_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3676),
            .ce(N__3398),
            .sr(_gnd_net_));
    defparam t0on_i14_LC_3_8_3.C_ON=1'b0;
    defparam t0on_i14_LC_3_8_3.SEQ_MODE=4'b1000;
    defparam t0on_i14_LC_3_8_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0on_i14_LC_3_8_3 (
            .in0(N__3297),
            .in1(N__3008),
            .in2(_gnd_net_),
            .in3(N__2975),
            .lcout(t0on_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3676),
            .ce(N__3398),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i12_1_lut_LC_3_8_4.C_ON=1'b0;
    defparam sub_34_inv_0_i12_1_lut_LC_3_8_4.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i12_1_lut_LC_3_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i12_1_lut_LC_3_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2956),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sub_34_inv_0_i10_1_lut_LC_3_8_5.C_ON=1'b0;
    defparam sub_34_inv_0_i10_1_lut_LC_3_8_5.SEQ_MODE=4'b0000;
    defparam sub_34_inv_0_i10_1_lut_LC_3_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 sub_34_inv_0_i10_1_lut_LC_3_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2917),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0off_i3_LC_3_9_0.C_ON=1'b0;
    defparam t0off_i3_LC_3_9_0.SEQ_MODE=4'b1000;
    defparam t0off_i3_LC_3_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i3_LC_3_9_0 (
            .in0(N__2879),
            .in1(N__3815),
            .in2(_gnd_net_),
            .in3(N__2870),
            .lcout(t0off_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i8_LC_3_9_1.C_ON=1'b0;
    defparam t0off_i8_LC_3_9_1.SEQ_MODE=4'b1000;
    defparam t0off_i8_LC_3_9_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0off_i8_LC_3_9_1 (
            .in0(N__3817),
            .in1(N__2864),
            .in2(_gnd_net_),
            .in3(N__2852),
            .lcout(t0off_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i2_LC_3_9_2.C_ON=1'b0;
    defparam t0off_i2_LC_3_9_2.SEQ_MODE=4'b1000;
    defparam t0off_i2_LC_3_9_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i2_LC_3_9_2 (
            .in0(N__2846),
            .in1(N__3814),
            .in2(_gnd_net_),
            .in3(N__2837),
            .lcout(t0off_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i10_LC_3_9_3.C_ON=1'b0;
    defparam t0off_i10_LC_3_9_3.SEQ_MODE=4'b1000;
    defparam t0off_i10_LC_3_9_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 t0off_i10_LC_3_9_3 (
            .in0(N__3812),
            .in1(_gnd_net_),
            .in2(N__2831),
            .in3(N__2816),
            .lcout(t0off_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i13_LC_3_9_4.C_ON=1'b0;
    defparam t0off_i13_LC_3_9_4.SEQ_MODE=4'b1000;
    defparam t0off_i13_LC_3_9_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i13_LC_3_9_4 (
            .in0(N__3161),
            .in1(N__3813),
            .in2(_gnd_net_),
            .in3(N__3149),
            .lcout(t0off_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i7_LC_3_9_7.C_ON=1'b0;
    defparam t0off_i7_LC_3_9_7.SEQ_MODE=4'b1000;
    defparam t0off_i7_LC_3_9_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0off_i7_LC_3_9_7 (
            .in0(N__3816),
            .in1(N__3143),
            .in2(_gnd_net_),
            .in3(N__3134),
            .lcout(t0off_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3677),
            .ce(N__3540),
            .sr(_gnd_net_));
    defparam t0off_i12_LC_3_10_1.C_ON=1'b0;
    defparam t0off_i12_LC_3_10_1.SEQ_MODE=4'b1000;
    defparam t0off_i12_LC_3_10_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i12_LC_3_10_1 (
            .in0(N__3128),
            .in1(N__3820),
            .in2(_gnd_net_),
            .in3(N__3119),
            .lcout(t0off_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam t0off_i9_LC_3_10_2.C_ON=1'b0;
    defparam t0off_i9_LC_3_10_2.SEQ_MODE=4'b1000;
    defparam t0off_i9_LC_3_10_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 t0off_i9_LC_3_10_2 (
            .in0(N__3824),
            .in1(N__3113),
            .in2(_gnd_net_),
            .in3(N__3107),
            .lcout(t0off_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam t0off_i14_LC_3_10_3.C_ON=1'b0;
    defparam t0off_i14_LC_3_10_3.SEQ_MODE=4'b1000;
    defparam t0off_i14_LC_3_10_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i14_LC_3_10_3 (
            .in0(N__3098),
            .in1(N__3821),
            .in2(_gnd_net_),
            .in3(N__3089),
            .lcout(t0off_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam t0off_i4_LC_3_10_4.C_ON=1'b0;
    defparam t0off_i4_LC_3_10_4.SEQ_MODE=4'b1000;
    defparam t0off_i4_LC_3_10_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0off_i4_LC_3_10_4 (
            .in0(N__3823),
            .in1(N__3083),
            .in2(_gnd_net_),
            .in3(N__3071),
            .lcout(t0off_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam t0off_i1_LC_3_10_5.C_ON=1'b0;
    defparam t0off_i1_LC_3_10_5.SEQ_MODE=4'b1000;
    defparam t0off_i1_LC_3_10_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i1_LC_3_10_5 (
            .in0(N__3065),
            .in1(N__3822),
            .in2(_gnd_net_),
            .in3(N__3053),
            .lcout(t0off_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam t0off_i0_LC_3_10_7.C_ON=1'b0;
    defparam t0off_i0_LC_3_10_7.SEQ_MODE=4'b1000;
    defparam t0off_i0_LC_3_10_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 t0off_i0_LC_3_10_7 (
            .in0(N__3047),
            .in1(N__3035),
            .in2(_gnd_net_),
            .in3(N__3819),
            .lcout(t0off_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3675),
            .ce(N__3541),
            .sr(_gnd_net_));
    defparam div_state_i1_LC_5_7_0.C_ON=1'b0;
    defparam div_state_i1_LC_5_7_0.SEQ_MODE=4'b1000;
    defparam div_state_i1_LC_5_7_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 div_state_i1_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__3277),
            .in2(_gnd_net_),
            .in3(N__3762),
            .lcout(div_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3692),
            .ce(N__3443),
            .sr(_gnd_net_));
    defparam i206_4_lut_LC_5_8_0.C_ON=1'b0;
    defparam i206_4_lut_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam i206_4_lut_LC_5_8_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i206_4_lut_LC_5_8_0 (
            .in0(N__3494),
            .in1(N__3482),
            .in2(N__3470),
            .in3(N__3458),
            .lcout(n441),
            .ltout(n441_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i214_2_lut_4_lut_LC_5_8_1.C_ON=1'b0;
    defparam i214_2_lut_4_lut_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam i214_2_lut_4_lut_LC_5_8_1.LUT_INIT=16'b0011011110111111;
    LogicCell40 i214_2_lut_4_lut_LC_5_8_1 (
            .in0(N__3757),
            .in1(N__3276),
            .in2(N__3446),
            .in3(N__3169),
            .lcout(n6_adj_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam div_state_i0_LC_5_8_3.C_ON=1'b0;
    defparam div_state_i0_LC_5_8_3.SEQ_MODE=4'b1000;
    defparam div_state_i0_LC_5_8_3.LUT_INIT=16'b1110111101001111;
    LogicCell40 div_state_i0_LC_5_8_3 (
            .in0(N__3758),
            .in1(N__3431),
            .in2(N__3293),
            .in3(N__3170),
            .lcout(div_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3689),
            .ce(),
            .sr(_gnd_net_));
    defparam i217_2_lut_LC_5_8_4.C_ON=1'b0;
    defparam i217_2_lut_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam i217_2_lut_LC_5_8_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 i217_2_lut_LC_5_8_4 (
            .in0(_gnd_net_),
            .in1(N__3271),
            .in2(_gnd_net_),
            .in3(N__3755),
            .lcout(n386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i218_1_lut_LC_5_8_5.C_ON=1'b0;
    defparam i218_1_lut_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam i218_1_lut_LC_5_8_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 i218_1_lut_LC_5_8_5 (
            .in0(N__3754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(div_state_1__N_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i208_2_lut_LC_5_8_6.C_ON=1'b0;
    defparam i208_2_lut_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam i208_2_lut_LC_5_8_6.LUT_INIT=16'b1100110000110011;
    LogicCell40 i208_2_lut_LC_5_8_6 (
            .in0(_gnd_net_),
            .in1(N__3272),
            .in2(_gnd_net_),
            .in3(N__3756),
            .lcout(n307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_5_9_1.C_ON=1'b0;
    defparam i11_4_lut_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_5_9_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_LC_5_9_1 (
            .in0(N__3239),
            .in1(N__3221),
            .in2(N__3206),
            .in3(N__3188),
            .lcout(),
            .ltout(n27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i205_4_lut_LC_5_9_2.C_ON=1'b0;
    defparam i205_4_lut_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam i205_4_lut_LC_5_9_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i205_4_lut_LC_5_9_2 (
            .in0(N__3971),
            .in1(N__4025),
            .in2(N__3173),
            .in3(N__3917),
            .lcout(n442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_5_9_4.C_ON=1'b0;
    defparam i10_4_lut_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_5_9_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_LC_5_9_4 (
            .in0(N__4072),
            .in1(N__4054),
            .in2(N__3889),
            .in3(N__4040),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_3_LC_5_10_0.C_ON=1'b0;
    defparam i12_4_lut_adj_3_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_3_LC_5_10_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_3_LC_5_10_0 (
            .in0(N__3703),
            .in1(N__4019),
            .in2(N__4004),
            .in3(N__3985),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i202_4_lut_LC_5_10_2.C_ON=1'b0;
    defparam i202_4_lut_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam i202_4_lut_LC_5_10_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 i202_4_lut_LC_5_10_2 (
            .in0(N__3847),
            .in1(N__3965),
            .in2(N__3950),
            .in3(N__3932),
            .lcout(n444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam t0off_i5_LC_6_9_0.C_ON=1'b0;
    defparam t0off_i5_LC_6_9_0.SEQ_MODE=4'b1000;
    defparam t0off_i5_LC_6_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i5_LC_6_9_0 (
            .in0(N__3911),
            .in1(N__3780),
            .in2(_gnd_net_),
            .in3(N__3902),
            .lcout(t0off_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3690),
            .ce(N__3529),
            .sr(_gnd_net_));
    defparam t0off_i6_LC_6_9_1.C_ON=1'b0;
    defparam t0off_i6_LC_6_9_1.SEQ_MODE=4'b1000;
    defparam t0off_i6_LC_6_9_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 t0off_i6_LC_6_9_1 (
            .in0(N__3781),
            .in1(N__3869),
            .in2(_gnd_net_),
            .in3(N__3860),
            .lcout(t0off_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3690),
            .ce(N__3529),
            .sr(_gnd_net_));
    defparam t0off_i11_LC_6_10_6.C_ON=1'b0;
    defparam t0off_i11_LC_6_10_6.SEQ_MODE=4'b1000;
    defparam t0off_i11_LC_6_10_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 t0off_i11_LC_6_10_6 (
            .in0(N__3836),
            .in1(N__3818),
            .in2(_gnd_net_),
            .in3(N__3716),
            .lcout(t0off_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3688),
            .ce(N__3533),
            .sr(_gnd_net_));
endmodule // vdc_gen_clk
